magic
tech scmos
timestamp 1701513645
<< nwell >>
rect 1540 298 1596 319
rect 1602 298 1632 319
rect 1683 297 1733 315
rect 1739 295 1768 316
rect 1827 299 1877 317
rect 1883 297 1912 318
rect 1970 300 2020 318
rect 2026 298 2055 319
rect 957 215 1014 233
rect 1020 213 1049 234
rect 1089 213 1118 234
rect 1124 215 1181 233
rect 1532 181 1588 202
rect 1770 184 1826 205
rect 2003 184 2059 205
rect 2241 187 2297 208
rect 1004 142 1025 171
rect 791 100 812 129
rect 794 44 811 93
rect 1007 86 1024 135
rect 1135 128 1156 157
rect 1332 148 1353 177
rect 1000 46 1021 75
rect 1138 72 1155 121
rect 1335 92 1352 141
rect 1441 131 1462 161
rect 787 4 808 33
rect 1131 32 1152 61
rect 1328 52 1349 81
rect 1441 69 1462 125
rect 1525 86 1546 142
rect 1573 86 1594 142
rect 1679 134 1700 164
rect 1531 53 1587 74
rect 1679 72 1700 128
rect 1763 89 1784 145
rect 1811 89 1832 145
rect 1912 134 1933 164
rect 1769 56 1825 77
rect 1912 72 1933 128
rect 1996 89 2017 145
rect 2044 89 2065 145
rect 2150 137 2171 167
rect 2002 56 2058 77
rect 2150 75 2171 131
rect 2234 92 2255 148
rect 2282 92 2303 148
rect 2370 130 2391 160
rect 2440 134 2470 155
rect 2486 134 2542 155
rect 2240 59 2296 80
rect 2370 58 2391 114
rect 847 -37 868 -8
rect 935 -32 956 -3
rect 1163 -23 1184 6
rect 1265 -25 1286 4
rect 1428 0 1449 30
rect 1666 3 1687 33
rect 1899 3 1920 33
rect 2137 6 2158 36
rect 2440 15 2470 36
rect 2486 15 2542 36
rect 850 -93 867 -44
rect 938 -88 955 -39
rect 1166 -79 1183 -30
rect 1268 -81 1285 -32
rect 1428 -90 1449 -34
rect 1532 -43 1588 -22
rect 843 -133 864 -104
rect 931 -128 952 -99
rect 1159 -119 1180 -90
rect 1261 -121 1282 -92
rect 1429 -141 1450 -111
rect 1525 -138 1546 -82
rect 1573 -138 1594 -82
rect 1666 -87 1687 -31
rect 1770 -40 1826 -19
rect 1667 -138 1688 -108
rect 1763 -135 1784 -79
rect 1811 -135 1832 -79
rect 1899 -87 1920 -31
rect 2003 -40 2059 -19
rect 1900 -138 1921 -108
rect 1996 -135 2017 -79
rect 2044 -135 2065 -79
rect 2137 -84 2158 -28
rect 2241 -37 2297 -16
rect 2370 -29 2391 1
rect 2440 -25 2470 -4
rect 2486 -25 2542 -4
rect 2138 -135 2159 -105
rect 2234 -132 2255 -76
rect 2282 -132 2303 -76
rect 2370 -101 2391 -45
rect 2440 -144 2470 -123
rect 2486 -144 2542 -123
rect 1000 -213 1021 -183
rect 1150 -213 1171 -183
rect 1297 -213 1318 -183
rect 1381 -196 1402 -166
rect 1531 -171 1587 -150
rect 1769 -168 1825 -147
rect 2002 -168 2058 -147
rect 2240 -165 2296 -144
rect 599 -285 616 -256
rect 599 -340 616 -291
rect 785 -305 806 -275
rect 941 -305 962 -275
rect 1000 -285 1021 -229
rect 1091 -305 1112 -275
rect 1150 -285 1171 -229
rect 1238 -305 1259 -275
rect 1297 -285 1318 -229
rect 1381 -268 1402 -212
rect 1429 -231 1450 -175
rect 1667 -228 1688 -172
rect 1900 -228 1921 -172
rect 2138 -225 2159 -169
rect 2369 -183 2390 -153
rect 2439 -179 2469 -158
rect 2485 -179 2541 -158
rect 1455 -275 1511 -254
rect 1693 -272 1749 -251
rect 1926 -272 1982 -251
rect 2164 -269 2220 -248
rect 2369 -255 2390 -199
rect 2439 -298 2469 -277
rect 2485 -298 2541 -277
rect 599 -398 616 -369
rect 661 -383 682 -327
rect 785 -333 841 -312
rect 941 -333 997 -312
rect 1091 -333 1147 -312
rect 1238 -333 1294 -312
rect 1448 -370 1469 -314
rect 1496 -370 1517 -314
rect 1686 -367 1707 -311
rect 1734 -367 1755 -311
rect 1919 -367 1940 -311
rect 1967 -367 1988 -311
rect 2157 -364 2178 -308
rect 2205 -364 2226 -308
rect 2369 -342 2390 -312
rect 2439 -338 2469 -317
rect 2485 -338 2541 -317
rect 599 -453 616 -404
rect 661 -419 682 -389
rect 778 -428 799 -372
rect 826 -428 847 -372
rect 934 -428 955 -372
rect 982 -428 1003 -372
rect 1084 -428 1105 -372
rect 1132 -428 1153 -372
rect 1231 -428 1252 -372
rect 1279 -428 1300 -372
rect 1454 -403 1510 -382
rect 1692 -400 1748 -379
rect 1925 -400 1981 -379
rect 2163 -397 2219 -376
rect 2369 -414 2390 -358
rect 784 -461 840 -440
rect 940 -461 996 -440
rect 1090 -461 1146 -440
rect 1237 -461 1293 -440
rect 2439 -457 2469 -436
rect 2485 -457 2541 -436
rect 459 -496 476 -467
rect 599 -506 616 -477
rect 599 -561 616 -512
rect 750 -536 771 -506
rect 863 -536 884 -506
rect 906 -536 927 -506
rect 1019 -536 1040 -506
rect 1056 -536 1077 -506
rect 1169 -536 1190 -506
rect 1212 -536 1233 -506
rect 1325 -536 1346 -506
rect 1458 -536 1479 -506
rect 1578 -536 1599 -506
rect 1697 -535 1718 -505
rect 1816 -535 1837 -505
rect 1930 -535 1951 -505
rect 2049 -535 2070 -505
rect 2151 -535 2172 -505
rect 2270 -535 2291 -505
rect 2352 -538 2373 -508
rect 457 -602 474 -573
rect 599 -617 616 -588
rect 750 -623 771 -567
rect 863 -623 884 -567
rect 906 -623 927 -567
rect 1019 -623 1040 -567
rect 1056 -623 1077 -567
rect 1169 -623 1190 -567
rect 1212 -623 1233 -567
rect 1325 -623 1346 -567
rect 1458 -613 1479 -557
rect 1578 -613 1599 -557
rect 1697 -612 1718 -556
rect 1816 -612 1837 -556
rect 1930 -612 1951 -556
rect 2049 -612 2070 -556
rect 2151 -612 2172 -556
rect 2270 -612 2291 -556
rect 2352 -615 2373 -559
rect 599 -672 616 -623
<< ntransistor >>
rect 1558 336 1561 344
rect 1575 336 1578 344
rect 1615 336 1618 344
rect 1695 338 1698 344
rect 1705 338 1708 344
rect 1715 338 1718 344
rect 1752 333 1755 341
rect 1839 340 1842 346
rect 1849 340 1852 346
rect 1859 340 1862 346
rect 1896 335 1899 343
rect 1982 341 1985 347
rect 1992 341 1995 347
rect 2002 341 2005 347
rect 2039 336 2042 344
rect 969 256 972 262
rect 979 256 982 262
rect 989 256 992 262
rect 999 256 1002 262
rect 1033 251 1036 259
rect 1102 251 1105 259
rect 1136 256 1139 262
rect 1146 256 1149 262
rect 1156 256 1159 262
rect 1166 256 1169 262
rect 1307 161 1315 164
rect 979 155 987 158
rect 1550 156 1553 164
rect 1567 156 1570 164
rect 1788 159 1791 167
rect 1805 159 1808 167
rect 2021 159 2024 167
rect 2038 159 2041 167
rect 2259 162 2262 170
rect 2276 162 2279 170
rect 1110 141 1118 144
rect 1479 144 1487 147
rect 1717 147 1725 150
rect 1950 147 1958 150
rect 2188 150 2196 153
rect 2408 143 2416 146
rect 1308 126 1313 129
rect 980 120 985 123
rect 766 113 774 116
rect 1500 121 1508 124
rect 1308 116 1313 119
rect 980 110 985 113
rect 1111 106 1116 109
rect 1308 106 1313 109
rect 980 100 985 103
rect 1738 124 1746 127
rect 1611 121 1619 124
rect 1479 104 1487 107
rect 1500 104 1508 107
rect 1111 96 1116 99
rect 1111 86 1116 89
rect 1611 104 1619 107
rect 1849 124 1857 127
rect 1971 124 1979 127
rect 1717 107 1725 110
rect 1738 107 1746 110
rect 1479 87 1487 90
rect 1849 107 1857 110
rect 2209 127 2217 130
rect 2082 124 2090 127
rect 1950 107 1958 110
rect 1971 107 1979 110
rect 1717 90 1725 93
rect 767 78 772 81
rect 2082 107 2090 110
rect 2320 127 2328 130
rect 2188 110 2196 113
rect 2209 110 2217 113
rect 1950 90 1958 93
rect 2320 110 2328 113
rect 2454 109 2457 117
rect 2504 109 2507 117
rect 2521 109 2524 117
rect 2188 93 2196 96
rect 2408 93 2416 96
rect 767 68 772 71
rect 2408 76 2416 79
rect 1303 65 1311 68
rect 767 58 772 61
rect 975 59 983 62
rect 1106 45 1114 48
rect 2454 53 2457 61
rect 2504 53 2507 61
rect 2521 53 2524 61
rect 1549 27 1552 35
rect 1566 27 1569 35
rect 1787 30 1790 38
rect 1804 30 1807 38
rect 2020 30 2023 38
rect 2037 30 2040 38
rect 2258 33 2261 41
rect 2275 33 2278 41
rect 762 17 770 20
rect 1466 13 1474 16
rect 1704 16 1712 19
rect 1937 16 1945 19
rect 2175 19 2183 22
rect 1138 -10 1146 -7
rect 822 -24 830 -21
rect 910 -19 918 -16
rect 1240 -12 1248 -9
rect 2408 -16 2416 -13
rect 1139 -45 1144 -42
rect 911 -54 916 -51
rect 823 -59 828 -56
rect 1241 -47 1246 -44
rect 1139 -55 1144 -52
rect 911 -64 916 -61
rect 1241 -57 1246 -54
rect 1466 -55 1474 -52
rect 823 -69 828 -66
rect 1139 -65 1144 -62
rect 911 -74 916 -71
rect 823 -79 828 -76
rect 1241 -67 1246 -64
rect 1704 -52 1712 -49
rect 1550 -68 1553 -60
rect 1567 -68 1570 -60
rect 1937 -52 1945 -49
rect 1788 -65 1791 -57
rect 1805 -65 1808 -57
rect 1466 -72 1474 -69
rect 1704 -69 1712 -66
rect 2175 -49 2183 -46
rect 2021 -65 2024 -57
rect 2038 -65 2041 -57
rect 2454 -50 2457 -42
rect 2504 -50 2507 -42
rect 2521 -50 2524 -42
rect 2259 -62 2262 -54
rect 2276 -62 2279 -54
rect 1937 -69 1945 -66
rect 2175 -66 2183 -63
rect 2408 -66 2416 -63
rect 2408 -83 2416 -80
rect 1134 -106 1142 -103
rect 818 -120 826 -117
rect 906 -115 914 -112
rect 1236 -108 1244 -105
rect 1500 -103 1508 -100
rect 1738 -100 1746 -97
rect 1611 -103 1619 -100
rect 1500 -120 1508 -117
rect 1467 -128 1475 -125
rect 1849 -100 1857 -97
rect 1971 -100 1979 -97
rect 1611 -120 1619 -117
rect 1738 -117 1746 -114
rect 1705 -125 1713 -122
rect 2209 -97 2217 -94
rect 2082 -100 2090 -97
rect 1849 -117 1857 -114
rect 1971 -117 1979 -114
rect 1938 -125 1946 -122
rect 2320 -97 2328 -94
rect 2082 -117 2090 -114
rect 2209 -114 2217 -111
rect 2176 -122 2184 -119
rect 2454 -106 2457 -98
rect 2504 -106 2507 -98
rect 2521 -106 2524 -98
rect 2320 -114 2328 -111
rect 1356 -183 1364 -180
rect 975 -200 983 -197
rect 1125 -200 1133 -197
rect 1272 -200 1280 -197
rect 1467 -196 1475 -193
rect 1549 -197 1552 -189
rect 1566 -197 1569 -189
rect 1705 -193 1713 -190
rect 1787 -194 1790 -186
rect 1804 -194 1807 -186
rect 1938 -193 1946 -190
rect 1467 -213 1475 -210
rect 1705 -210 1713 -207
rect 2020 -194 2023 -186
rect 2037 -194 2040 -186
rect 2407 -170 2415 -167
rect 2176 -190 2184 -187
rect 2258 -191 2261 -183
rect 2275 -191 2278 -183
rect 1938 -210 1946 -207
rect 2176 -207 2184 -204
rect 2453 -204 2456 -196
rect 2503 -204 2506 -196
rect 2520 -204 2523 -196
rect 2407 -220 2415 -217
rect 1356 -233 1364 -230
rect 975 -250 983 -247
rect 572 -272 577 -269
rect 1125 -250 1133 -247
rect 975 -267 983 -264
rect 1272 -250 1280 -247
rect 1125 -267 1133 -264
rect 2407 -237 2415 -234
rect 1356 -250 1364 -247
rect 1272 -267 1280 -264
rect 2453 -260 2456 -252
rect 2503 -260 2506 -252
rect 2520 -260 2523 -252
rect 760 -292 768 -289
rect 916 -292 924 -289
rect 1066 -292 1074 -289
rect 1213 -292 1221 -289
rect 1473 -300 1476 -292
rect 1490 -300 1493 -292
rect 1711 -297 1714 -289
rect 1728 -297 1731 -289
rect 1944 -297 1947 -289
rect 1961 -297 1964 -289
rect 2182 -294 2185 -286
rect 2199 -294 2202 -286
rect 572 -306 577 -303
rect 572 -316 577 -313
rect 572 -326 577 -323
rect 699 -348 707 -345
rect 1423 -335 1431 -332
rect 1661 -332 1669 -329
rect 1534 -335 1542 -332
rect 803 -358 806 -350
rect 820 -358 823 -350
rect 959 -358 962 -350
rect 976 -358 979 -350
rect 1109 -358 1112 -350
rect 1126 -358 1129 -350
rect 1256 -358 1259 -350
rect 1273 -358 1276 -350
rect 1423 -352 1431 -349
rect 1772 -332 1780 -329
rect 1894 -332 1902 -329
rect 1661 -349 1669 -346
rect 1534 -352 1542 -349
rect 2132 -329 2140 -326
rect 2005 -332 2013 -329
rect 1772 -349 1780 -346
rect 1894 -349 1902 -346
rect 2243 -329 2251 -326
rect 2132 -346 2140 -343
rect 2005 -349 2013 -346
rect 2407 -329 2415 -326
rect 2243 -346 2251 -343
rect 699 -365 707 -362
rect 2453 -363 2456 -355
rect 2503 -363 2506 -355
rect 2520 -363 2523 -355
rect 2407 -379 2415 -376
rect 572 -385 577 -382
rect 753 -393 761 -390
rect 699 -405 707 -402
rect 864 -393 872 -390
rect 909 -393 917 -390
rect 753 -410 761 -407
rect 572 -419 577 -416
rect 1020 -393 1028 -390
rect 1059 -393 1067 -390
rect 864 -410 872 -407
rect 909 -410 917 -407
rect 1170 -393 1178 -390
rect 1206 -393 1214 -390
rect 1020 -410 1028 -407
rect 1059 -410 1067 -407
rect 1317 -393 1325 -390
rect 1170 -410 1178 -407
rect 1206 -410 1214 -407
rect 1317 -410 1325 -407
rect 2407 -396 2415 -393
rect 572 -429 577 -426
rect 1472 -429 1475 -421
rect 1489 -429 1492 -421
rect 1710 -426 1713 -418
rect 1727 -426 1730 -418
rect 1943 -426 1946 -418
rect 1960 -426 1963 -418
rect 2181 -423 2184 -415
rect 2198 -423 2201 -415
rect 2453 -419 2456 -411
rect 2503 -419 2506 -411
rect 2520 -419 2523 -411
rect 572 -439 577 -436
rect 498 -483 503 -480
rect 802 -487 805 -479
rect 819 -487 822 -479
rect 958 -487 961 -479
rect 975 -487 978 -479
rect 1108 -487 1111 -479
rect 1125 -487 1128 -479
rect 1255 -487 1258 -479
rect 1272 -487 1275 -479
rect 572 -493 577 -490
rect 572 -527 577 -524
rect 788 -523 796 -520
rect 838 -523 846 -520
rect 944 -523 952 -520
rect 994 -523 1002 -520
rect 1094 -523 1102 -520
rect 1144 -523 1152 -520
rect 1250 -523 1258 -520
rect 1300 -523 1308 -520
rect 1496 -523 1504 -520
rect 1553 -523 1561 -520
rect 1735 -522 1743 -519
rect 1791 -522 1799 -519
rect 1968 -522 1976 -519
rect 2024 -522 2032 -519
rect 2189 -522 2197 -519
rect 2245 -522 2253 -519
rect 2327 -525 2335 -522
rect 572 -537 577 -534
rect 572 -547 577 -544
rect 1496 -578 1504 -575
rect 430 -589 435 -586
rect 788 -588 796 -585
rect 572 -604 577 -601
rect 838 -588 846 -585
rect 944 -588 952 -585
rect 788 -605 796 -602
rect 994 -588 1002 -585
rect 1094 -588 1102 -585
rect 838 -605 846 -602
rect 944 -605 952 -602
rect 1144 -588 1152 -585
rect 1250 -588 1258 -585
rect 994 -605 1002 -602
rect 1094 -605 1102 -602
rect 1300 -588 1308 -585
rect 1144 -605 1152 -602
rect 1250 -605 1258 -602
rect 1553 -578 1561 -575
rect 1735 -577 1743 -574
rect 1496 -595 1504 -592
rect 1300 -605 1308 -602
rect 1791 -577 1799 -574
rect 1968 -577 1976 -574
rect 1553 -595 1561 -592
rect 1735 -594 1743 -591
rect 2024 -577 2032 -574
rect 2189 -577 2197 -574
rect 1791 -594 1799 -591
rect 1968 -594 1976 -591
rect 2245 -577 2253 -574
rect 2024 -594 2032 -591
rect 2189 -594 2197 -591
rect 2327 -580 2335 -577
rect 2245 -594 2253 -591
rect 2327 -597 2335 -594
rect 572 -638 577 -635
rect 572 -648 577 -645
rect 572 -658 577 -655
<< ptransistor >>
rect 1558 304 1561 312
rect 1575 304 1578 312
rect 1615 304 1618 312
rect 1695 303 1698 309
rect 1705 303 1708 309
rect 1715 303 1718 309
rect 1752 301 1755 309
rect 1839 305 1842 311
rect 1849 305 1852 311
rect 1859 305 1862 311
rect 1896 303 1899 311
rect 1982 306 1985 312
rect 1992 306 1995 312
rect 2002 306 2005 312
rect 2039 304 2042 312
rect 969 221 972 227
rect 979 221 982 227
rect 989 221 992 227
rect 999 221 1002 227
rect 1033 219 1036 227
rect 1102 219 1105 227
rect 1136 221 1139 227
rect 1146 221 1149 227
rect 1156 221 1159 227
rect 1166 221 1169 227
rect 1550 188 1553 196
rect 1567 188 1570 196
rect 1788 191 1791 199
rect 1805 191 1808 199
rect 2021 191 2024 199
rect 2038 191 2041 199
rect 2259 194 2262 202
rect 2276 194 2279 202
rect 1339 161 1347 164
rect 1011 155 1019 158
rect 1447 144 1455 147
rect 1142 141 1150 144
rect 1685 147 1693 150
rect 1918 147 1926 150
rect 2156 150 2164 153
rect 2376 143 2384 146
rect 1341 126 1346 129
rect 1013 120 1018 123
rect 798 113 806 116
rect 1341 116 1346 119
rect 1013 110 1018 113
rect 1144 106 1149 109
rect 1013 100 1018 103
rect 1341 106 1346 109
rect 1532 121 1540 124
rect 1579 121 1587 124
rect 1447 104 1455 107
rect 1532 104 1540 107
rect 1144 96 1149 99
rect 1144 86 1149 89
rect 1579 104 1587 107
rect 1770 124 1778 127
rect 1817 124 1825 127
rect 1685 107 1693 110
rect 1770 107 1778 110
rect 1447 87 1455 90
rect 1817 107 1825 110
rect 2003 124 2011 127
rect 2050 124 2058 127
rect 1918 107 1926 110
rect 2003 107 2011 110
rect 1685 90 1693 93
rect 800 78 805 81
rect 2050 107 2058 110
rect 2454 141 2457 149
rect 2504 141 2507 149
rect 2521 141 2524 149
rect 2241 127 2249 130
rect 2288 127 2296 130
rect 2156 110 2164 113
rect 2241 110 2249 113
rect 1918 90 1926 93
rect 2288 110 2296 113
rect 2156 93 2164 96
rect 2376 93 2384 96
rect 800 68 805 71
rect 2376 76 2384 79
rect 800 58 805 61
rect 1335 65 1343 68
rect 1007 59 1015 62
rect 1549 60 1552 68
rect 1566 60 1569 68
rect 1787 63 1790 71
rect 1804 63 1807 71
rect 2020 63 2023 71
rect 2037 63 2040 71
rect 2258 66 2261 74
rect 2275 66 2278 74
rect 1138 45 1146 48
rect 794 17 802 20
rect 1434 13 1442 16
rect 1672 16 1680 19
rect 1905 16 1913 19
rect 2143 19 2151 22
rect 2454 21 2457 29
rect 2504 21 2507 29
rect 2521 21 2524 29
rect 854 -24 862 -21
rect 1170 -10 1178 -7
rect 942 -19 950 -16
rect 1272 -12 1280 -9
rect 2376 -16 2384 -13
rect 1550 -36 1553 -28
rect 1567 -36 1570 -28
rect 1788 -33 1791 -25
rect 1805 -33 1808 -25
rect 2021 -33 2024 -25
rect 2038 -33 2041 -25
rect 2259 -30 2262 -22
rect 2276 -30 2279 -22
rect 2454 -18 2457 -10
rect 2504 -18 2507 -10
rect 2521 -18 2524 -10
rect 1172 -45 1177 -42
rect 944 -54 949 -51
rect 856 -59 861 -56
rect 1274 -47 1279 -44
rect 1172 -55 1177 -52
rect 944 -64 949 -61
rect 1274 -57 1279 -54
rect 1434 -55 1442 -52
rect 856 -69 861 -66
rect 1172 -65 1177 -62
rect 1274 -67 1279 -64
rect 944 -74 949 -71
rect 1672 -52 1680 -49
rect 1905 -52 1913 -49
rect 1434 -72 1442 -69
rect 856 -79 861 -76
rect 1672 -69 1680 -66
rect 2143 -49 2151 -46
rect 1905 -69 1913 -66
rect 2143 -66 2151 -63
rect 2376 -66 2384 -63
rect 2376 -83 2384 -80
rect 850 -120 858 -117
rect 1166 -106 1174 -103
rect 938 -115 946 -112
rect 1268 -108 1276 -105
rect 1532 -103 1540 -100
rect 1579 -103 1587 -100
rect 1532 -120 1540 -117
rect 1435 -128 1443 -125
rect 1770 -100 1778 -97
rect 1817 -100 1825 -97
rect 1579 -120 1587 -117
rect 1770 -117 1778 -114
rect 1673 -125 1681 -122
rect 2003 -100 2011 -97
rect 2050 -100 2058 -97
rect 1817 -117 1825 -114
rect 2003 -117 2011 -114
rect 1906 -125 1914 -122
rect 2241 -97 2249 -94
rect 2288 -97 2296 -94
rect 2050 -117 2058 -114
rect 2241 -114 2249 -111
rect 2144 -122 2152 -119
rect 2288 -114 2296 -111
rect 2454 -138 2457 -130
rect 2504 -138 2507 -130
rect 2521 -138 2524 -130
rect 1549 -164 1552 -156
rect 1566 -164 1569 -156
rect 1787 -161 1790 -153
rect 1804 -161 1807 -153
rect 2020 -161 2023 -153
rect 2037 -161 2040 -153
rect 2258 -158 2261 -150
rect 2275 -158 2278 -150
rect 1388 -183 1396 -180
rect 1007 -200 1015 -197
rect 1157 -200 1165 -197
rect 1435 -196 1443 -193
rect 1304 -200 1312 -197
rect 1673 -193 1681 -190
rect 1906 -193 1914 -190
rect 1435 -213 1443 -210
rect 1673 -210 1681 -207
rect 2375 -170 2383 -167
rect 2453 -172 2456 -164
rect 2503 -172 2506 -164
rect 2520 -172 2523 -164
rect 2144 -190 2152 -187
rect 1906 -210 1914 -207
rect 2144 -207 2152 -204
rect 2375 -220 2383 -217
rect 1388 -233 1396 -230
rect 1007 -250 1015 -247
rect 1157 -250 1165 -247
rect 1007 -267 1015 -264
rect 605 -272 610 -269
rect 1304 -250 1312 -247
rect 1157 -267 1165 -264
rect 2375 -237 2383 -234
rect 1388 -250 1396 -247
rect 1304 -267 1312 -264
rect 1473 -268 1476 -260
rect 1490 -268 1493 -260
rect 1711 -265 1714 -257
rect 1728 -265 1731 -257
rect 1944 -265 1947 -257
rect 1961 -265 1964 -257
rect 2182 -262 2185 -254
rect 2199 -262 2202 -254
rect 792 -292 800 -289
rect 948 -292 956 -289
rect 1098 -292 1106 -289
rect 1245 -292 1253 -289
rect 2453 -292 2456 -284
rect 2503 -292 2506 -284
rect 2520 -292 2523 -284
rect 605 -306 610 -303
rect 605 -316 610 -313
rect 605 -326 610 -323
rect 803 -326 806 -318
rect 820 -326 823 -318
rect 959 -326 962 -318
rect 976 -326 979 -318
rect 1109 -326 1112 -318
rect 1126 -326 1129 -318
rect 1256 -326 1259 -318
rect 1273 -326 1276 -318
rect 667 -348 675 -345
rect 1455 -335 1463 -332
rect 1502 -335 1510 -332
rect 1455 -352 1463 -349
rect 1693 -332 1701 -329
rect 1740 -332 1748 -329
rect 1693 -349 1701 -346
rect 1502 -352 1510 -349
rect 1926 -332 1934 -329
rect 1973 -332 1981 -329
rect 1740 -349 1748 -346
rect 1926 -349 1934 -346
rect 2164 -329 2172 -326
rect 2211 -329 2219 -326
rect 2375 -329 2383 -326
rect 2164 -346 2172 -343
rect 1973 -349 1981 -346
rect 2453 -331 2456 -323
rect 2503 -331 2506 -323
rect 2520 -331 2523 -323
rect 2211 -346 2219 -343
rect 667 -365 675 -362
rect 2375 -379 2383 -376
rect 605 -385 610 -382
rect 667 -405 675 -402
rect 785 -393 793 -390
rect 832 -393 840 -390
rect 785 -410 793 -407
rect 605 -419 610 -416
rect 941 -393 949 -390
rect 988 -393 996 -390
rect 832 -410 840 -407
rect 941 -410 949 -407
rect 1091 -393 1099 -390
rect 1138 -393 1146 -390
rect 988 -410 996 -407
rect 1091 -410 1099 -407
rect 1238 -393 1246 -390
rect 1285 -393 1293 -390
rect 1138 -410 1146 -407
rect 1238 -410 1246 -407
rect 1472 -396 1475 -388
rect 1489 -396 1492 -388
rect 1710 -393 1713 -385
rect 1727 -393 1730 -385
rect 1943 -393 1946 -385
rect 1960 -393 1963 -385
rect 2181 -390 2184 -382
rect 2198 -390 2201 -382
rect 1285 -410 1293 -407
rect 2375 -396 2383 -393
rect 605 -429 610 -426
rect 605 -439 610 -436
rect 802 -454 805 -446
rect 819 -454 822 -446
rect 958 -454 961 -446
rect 975 -454 978 -446
rect 1108 -454 1111 -446
rect 1125 -454 1128 -446
rect 1255 -454 1258 -446
rect 1272 -454 1275 -446
rect 2453 -451 2456 -443
rect 2503 -451 2506 -443
rect 2520 -451 2523 -443
rect 465 -483 470 -480
rect 605 -493 610 -490
rect 756 -523 764 -520
rect 605 -527 610 -524
rect 870 -523 878 -520
rect 912 -523 920 -520
rect 1026 -523 1034 -520
rect 1062 -523 1070 -520
rect 1176 -523 1184 -520
rect 1218 -523 1226 -520
rect 1332 -523 1340 -520
rect 1464 -523 1472 -520
rect 1585 -523 1593 -520
rect 1703 -522 1711 -519
rect 1823 -522 1831 -519
rect 1936 -522 1944 -519
rect 2056 -522 2064 -519
rect 2157 -522 2165 -519
rect 2277 -522 2285 -519
rect 2359 -525 2367 -522
rect 605 -537 610 -534
rect 605 -547 610 -544
rect 1464 -578 1472 -575
rect 463 -589 468 -586
rect 756 -588 764 -585
rect 605 -604 610 -601
rect 870 -588 878 -585
rect 912 -588 920 -585
rect 756 -605 764 -602
rect 1026 -588 1034 -585
rect 1062 -588 1070 -585
rect 870 -605 878 -602
rect 912 -605 920 -602
rect 1176 -588 1184 -585
rect 1218 -588 1226 -585
rect 1026 -605 1034 -602
rect 1062 -605 1070 -602
rect 1332 -588 1340 -585
rect 1176 -605 1184 -602
rect 1218 -605 1226 -602
rect 1585 -578 1593 -575
rect 1703 -577 1711 -574
rect 1464 -595 1472 -592
rect 1332 -605 1340 -602
rect 1823 -577 1831 -574
rect 1936 -577 1944 -574
rect 1585 -595 1593 -592
rect 1703 -594 1711 -591
rect 2056 -577 2064 -574
rect 2157 -577 2165 -574
rect 1823 -594 1831 -591
rect 1936 -594 1944 -591
rect 2277 -577 2285 -574
rect 2056 -594 2064 -591
rect 2157 -594 2165 -591
rect 2359 -580 2367 -577
rect 2277 -594 2285 -591
rect 2359 -597 2367 -594
rect 605 -638 610 -635
rect 605 -648 610 -645
rect 605 -658 610 -655
<< ndiffusion >>
rect 1554 336 1558 344
rect 1561 336 1565 344
rect 1570 336 1575 344
rect 1578 336 1581 344
rect 1612 336 1615 344
rect 1618 336 1622 344
rect 1694 338 1695 344
rect 1698 338 1699 344
rect 1704 338 1705 344
rect 1708 338 1709 344
rect 1714 338 1715 344
rect 1718 338 1719 344
rect 1724 338 1725 344
rect 1749 333 1752 341
rect 1755 333 1758 341
rect 1838 340 1839 346
rect 1842 340 1843 346
rect 1848 340 1849 346
rect 1852 340 1853 346
rect 1858 340 1859 346
rect 1862 340 1863 346
rect 1868 340 1869 346
rect 1893 335 1896 343
rect 1899 335 1902 343
rect 1981 341 1982 347
rect 1985 341 1986 347
rect 1991 341 1992 347
rect 1995 341 1996 347
rect 2001 341 2002 347
rect 2005 341 2006 347
rect 2011 341 2012 347
rect 2036 336 2039 344
rect 2042 336 2045 344
rect 968 256 969 262
rect 972 256 973 262
rect 978 256 979 262
rect 982 256 983 262
rect 988 256 989 262
rect 992 256 993 262
rect 998 256 999 262
rect 1002 256 1003 262
rect 1030 251 1033 259
rect 1036 251 1039 259
rect 1099 251 1102 259
rect 1105 251 1108 259
rect 1135 256 1136 262
rect 1139 256 1140 262
rect 1145 256 1146 262
rect 1149 256 1150 262
rect 1155 256 1156 262
rect 1159 256 1160 262
rect 1165 256 1166 262
rect 1169 256 1170 262
rect 979 158 987 161
rect 1307 164 1315 167
rect 979 152 987 155
rect 1307 158 1315 161
rect 1547 156 1550 164
rect 1553 156 1567 164
rect 1570 156 1578 164
rect 1785 159 1788 167
rect 1791 159 1805 167
rect 1808 159 1816 167
rect 2018 159 2021 167
rect 2024 159 2038 167
rect 2041 159 2049 167
rect 2256 162 2259 170
rect 2262 162 2276 170
rect 2279 162 2287 170
rect 1110 144 1118 147
rect 1110 138 1118 141
rect 1479 147 1487 151
rect 1717 150 1725 154
rect 1479 141 1487 144
rect 1717 144 1725 147
rect 1950 150 1958 154
rect 2188 153 2196 157
rect 1950 144 1958 147
rect 2188 147 2196 150
rect 2408 146 2416 150
rect 766 116 774 119
rect 980 123 985 124
rect 1308 129 1313 130
rect 766 110 774 113
rect 980 113 985 120
rect 1308 119 1313 126
rect 1500 124 1508 127
rect 980 103 985 110
rect 1111 109 1116 110
rect 1308 109 1313 116
rect 980 99 985 100
rect 1111 99 1116 106
rect 1308 105 1313 106
rect 1479 107 1487 110
rect 1500 107 1508 121
rect 1738 127 1746 130
rect 1611 124 1619 127
rect 1111 89 1116 96
rect 767 81 772 82
rect 1111 85 1116 86
rect 1479 99 1487 104
rect 1500 100 1508 104
rect 1611 107 1619 121
rect 1717 110 1725 113
rect 1738 110 1746 124
rect 1849 127 1857 130
rect 1971 127 1979 130
rect 1611 100 1619 104
rect 1479 90 1487 94
rect 1717 102 1725 107
rect 1738 103 1746 107
rect 1849 110 1857 124
rect 1849 103 1857 107
rect 1950 110 1958 113
rect 1971 110 1979 124
rect 2209 130 2217 133
rect 2082 127 2090 130
rect 1717 93 1725 97
rect 1479 83 1487 87
rect 1717 86 1725 90
rect 1950 102 1958 107
rect 1971 103 1979 107
rect 2082 110 2090 124
rect 2188 113 2196 116
rect 2209 113 2217 127
rect 2408 140 2416 143
rect 2320 130 2328 133
rect 2082 103 2090 107
rect 1950 93 1958 97
rect 2188 105 2196 110
rect 2209 106 2217 110
rect 2320 113 2328 127
rect 2320 106 2328 110
rect 2450 109 2454 117
rect 2457 109 2460 117
rect 2501 109 2504 117
rect 2507 109 2521 117
rect 2524 109 2528 117
rect 2188 96 2196 100
rect 2408 96 2416 99
rect 1950 86 1958 90
rect 2188 89 2196 93
rect 2408 79 2416 93
rect 767 71 772 78
rect 767 61 772 68
rect 975 62 983 65
rect 1303 68 1311 71
rect 767 57 772 58
rect 975 56 983 59
rect 1303 62 1311 65
rect 2408 72 2416 76
rect 1106 48 1114 51
rect 1106 42 1114 45
rect 2450 53 2454 61
rect 2457 53 2460 61
rect 2501 53 2504 61
rect 2507 53 2521 61
rect 2524 53 2528 61
rect 1545 27 1549 35
rect 1552 27 1566 35
rect 1569 27 1572 35
rect 1783 30 1787 38
rect 1790 30 1804 38
rect 1807 30 1810 38
rect 2016 30 2020 38
rect 2023 30 2037 38
rect 2040 30 2043 38
rect 2254 33 2258 41
rect 2261 33 2275 41
rect 2278 33 2281 41
rect 762 20 770 23
rect 762 14 770 17
rect 1466 16 1474 20
rect 1704 19 1712 23
rect 1466 10 1474 13
rect 1704 13 1712 16
rect 1937 19 1945 23
rect 2175 22 2183 26
rect 1937 13 1945 16
rect 2175 16 2183 19
rect 1138 -7 1146 -4
rect 822 -21 830 -18
rect 910 -16 918 -13
rect 822 -27 830 -24
rect 910 -22 918 -19
rect 1138 -13 1146 -10
rect 1240 -9 1248 -6
rect 1240 -15 1248 -12
rect 2408 -13 2416 -9
rect 2408 -19 2416 -16
rect 1139 -42 1144 -41
rect 823 -56 828 -55
rect 911 -51 916 -50
rect 823 -66 828 -59
rect 911 -61 916 -54
rect 1139 -52 1144 -45
rect 1241 -44 1246 -43
rect 1139 -62 1144 -55
rect 1241 -54 1246 -47
rect 1466 -52 1474 -49
rect 823 -76 828 -69
rect 911 -71 916 -64
rect 823 -80 828 -79
rect 911 -75 916 -74
rect 1139 -66 1144 -65
rect 1241 -64 1246 -57
rect 1241 -68 1246 -67
rect 1466 -69 1474 -55
rect 1704 -49 1712 -46
rect 1547 -68 1550 -60
rect 1553 -68 1567 -60
rect 1570 -68 1578 -60
rect 1704 -66 1712 -52
rect 1937 -49 1945 -46
rect 1785 -65 1788 -57
rect 1791 -65 1805 -57
rect 1808 -65 1816 -57
rect 1466 -76 1474 -72
rect 1704 -73 1712 -69
rect 1937 -66 1945 -52
rect 2175 -46 2183 -43
rect 2018 -65 2021 -57
rect 2024 -65 2038 -57
rect 2041 -65 2049 -57
rect 2175 -63 2183 -49
rect 2450 -50 2454 -42
rect 2457 -50 2460 -42
rect 2501 -50 2504 -42
rect 2507 -50 2521 -42
rect 2524 -50 2528 -42
rect 2256 -62 2259 -54
rect 2262 -62 2276 -54
rect 2279 -62 2287 -54
rect 1937 -73 1945 -69
rect 2175 -70 2183 -66
rect 2408 -63 2416 -60
rect 2408 -80 2416 -66
rect 1134 -103 1142 -100
rect 818 -117 826 -114
rect 906 -112 914 -109
rect 818 -123 826 -120
rect 906 -118 914 -115
rect 1134 -109 1142 -106
rect 1236 -105 1244 -102
rect 1500 -100 1508 -97
rect 1236 -111 1244 -108
rect 1500 -117 1508 -103
rect 1738 -97 1746 -94
rect 1611 -100 1619 -97
rect 1467 -125 1475 -121
rect 1500 -124 1508 -120
rect 1611 -117 1619 -103
rect 1738 -114 1746 -100
rect 1849 -97 1857 -94
rect 1971 -97 1979 -94
rect 1611 -124 1619 -120
rect 1705 -122 1713 -118
rect 1738 -121 1746 -117
rect 1849 -114 1857 -100
rect 1971 -114 1979 -100
rect 2209 -94 2217 -91
rect 2082 -97 2090 -94
rect 1849 -121 1857 -117
rect 1467 -131 1475 -128
rect 1705 -128 1713 -125
rect 1938 -122 1946 -118
rect 1971 -121 1979 -117
rect 2082 -114 2090 -100
rect 2209 -111 2217 -97
rect 2408 -87 2416 -83
rect 2320 -94 2328 -91
rect 2082 -121 2090 -117
rect 2176 -119 2184 -115
rect 2209 -118 2217 -114
rect 2320 -111 2328 -97
rect 2450 -106 2454 -98
rect 2457 -106 2460 -98
rect 2501 -106 2504 -98
rect 2507 -106 2521 -98
rect 2524 -106 2528 -98
rect 2320 -118 2328 -114
rect 1938 -128 1946 -125
rect 2176 -125 2184 -122
rect 1356 -180 1364 -176
rect 1356 -186 1364 -183
rect 975 -197 983 -193
rect 975 -203 983 -200
rect 1125 -197 1133 -193
rect 1125 -203 1133 -200
rect 1272 -197 1280 -193
rect 1467 -193 1475 -190
rect 1272 -203 1280 -200
rect 1467 -210 1475 -196
rect 1545 -197 1549 -189
rect 1552 -197 1566 -189
rect 1569 -197 1572 -189
rect 1705 -190 1713 -187
rect 1705 -207 1713 -193
rect 1783 -194 1787 -186
rect 1790 -194 1804 -186
rect 1807 -194 1810 -186
rect 1938 -190 1946 -187
rect 1467 -217 1475 -213
rect 1705 -214 1713 -210
rect 1938 -207 1946 -193
rect 2016 -194 2020 -186
rect 2023 -194 2037 -186
rect 2040 -194 2043 -186
rect 2407 -167 2415 -163
rect 2407 -173 2415 -170
rect 2176 -187 2184 -184
rect 2176 -204 2184 -190
rect 2254 -191 2258 -183
rect 2261 -191 2275 -183
rect 2278 -191 2281 -183
rect 1938 -214 1946 -210
rect 2176 -211 2184 -207
rect 2449 -204 2453 -196
rect 2456 -204 2459 -196
rect 2500 -204 2503 -196
rect 2506 -204 2520 -196
rect 2523 -204 2527 -196
rect 2407 -217 2415 -214
rect 1356 -230 1364 -227
rect 975 -247 983 -244
rect 572 -269 577 -266
rect 572 -275 577 -272
rect 975 -264 983 -250
rect 1125 -247 1133 -244
rect 975 -271 983 -267
rect 1125 -264 1133 -250
rect 1272 -247 1280 -244
rect 1125 -271 1133 -267
rect 1272 -264 1280 -250
rect 1356 -247 1364 -233
rect 2407 -234 2415 -220
rect 2407 -241 2415 -237
rect 1356 -254 1364 -250
rect 1272 -271 1280 -267
rect 2449 -260 2453 -252
rect 2456 -260 2459 -252
rect 2500 -260 2503 -252
rect 2506 -260 2520 -252
rect 2523 -260 2527 -252
rect 760 -289 768 -285
rect 760 -295 768 -292
rect 916 -289 924 -285
rect 572 -303 577 -301
rect 916 -295 924 -292
rect 1066 -289 1074 -285
rect 1066 -295 1074 -292
rect 1213 -289 1221 -285
rect 1213 -295 1221 -292
rect 1470 -300 1473 -292
rect 1476 -300 1490 -292
rect 1493 -300 1501 -292
rect 1708 -297 1711 -289
rect 1714 -297 1728 -289
rect 1731 -297 1739 -289
rect 1941 -297 1944 -289
rect 1947 -297 1961 -289
rect 1964 -297 1972 -289
rect 2179 -294 2182 -286
rect 2185 -294 2199 -286
rect 2202 -294 2210 -286
rect 572 -313 577 -306
rect 572 -323 577 -316
rect 572 -327 577 -326
rect 699 -345 707 -341
rect 699 -352 707 -348
rect 1423 -332 1431 -329
rect 1423 -349 1431 -335
rect 1661 -329 1669 -326
rect 1534 -332 1542 -329
rect 699 -362 707 -357
rect 800 -358 803 -350
rect 806 -358 820 -350
rect 823 -358 831 -350
rect 956 -358 959 -350
rect 962 -358 976 -350
rect 979 -358 987 -350
rect 1106 -358 1109 -350
rect 1112 -358 1126 -350
rect 1129 -358 1137 -350
rect 1253 -358 1256 -350
rect 1259 -358 1273 -350
rect 1276 -358 1284 -350
rect 1423 -356 1431 -352
rect 1534 -349 1542 -335
rect 1661 -346 1669 -332
rect 1772 -329 1780 -326
rect 1894 -329 1902 -326
rect 1534 -356 1542 -352
rect 1661 -353 1669 -349
rect 1772 -346 1780 -332
rect 1894 -346 1902 -332
rect 2132 -326 2140 -323
rect 2005 -329 2013 -326
rect 1772 -353 1780 -349
rect 1894 -353 1902 -349
rect 2005 -346 2013 -332
rect 2132 -343 2140 -329
rect 2243 -326 2251 -323
rect 2005 -353 2013 -349
rect 2132 -350 2140 -346
rect 2243 -343 2251 -329
rect 2407 -326 2415 -322
rect 2407 -332 2415 -329
rect 2243 -350 2251 -346
rect 2449 -363 2453 -355
rect 2456 -363 2459 -355
rect 2500 -363 2503 -355
rect 2506 -363 2520 -355
rect 2523 -363 2527 -355
rect 699 -368 707 -365
rect 572 -382 577 -379
rect 2407 -376 2415 -373
rect 572 -388 577 -385
rect 753 -390 761 -387
rect 699 -402 707 -399
rect 572 -416 577 -414
rect 699 -409 707 -405
rect 753 -407 761 -393
rect 864 -390 872 -387
rect 909 -390 917 -387
rect 753 -414 761 -410
rect 864 -407 872 -393
rect 909 -407 917 -393
rect 1020 -390 1028 -387
rect 1059 -390 1067 -387
rect 864 -414 872 -410
rect 909 -414 917 -410
rect 1020 -407 1028 -393
rect 1059 -407 1067 -393
rect 1170 -390 1178 -387
rect 1206 -390 1214 -387
rect 1020 -414 1028 -410
rect 1059 -414 1067 -410
rect 1170 -407 1178 -393
rect 1206 -407 1214 -393
rect 1317 -390 1325 -387
rect 1170 -414 1178 -410
rect 1206 -414 1214 -410
rect 1317 -407 1325 -393
rect 1317 -414 1325 -410
rect 572 -426 577 -419
rect 2407 -393 2415 -379
rect 2407 -400 2415 -396
rect 1468 -429 1472 -421
rect 1475 -429 1489 -421
rect 1492 -429 1495 -421
rect 1706 -426 1710 -418
rect 1713 -426 1727 -418
rect 1730 -426 1733 -418
rect 1939 -426 1943 -418
rect 1946 -426 1960 -418
rect 1963 -426 1966 -418
rect 2177 -423 2181 -415
rect 2184 -423 2198 -415
rect 2201 -423 2204 -415
rect 2449 -419 2453 -411
rect 2456 -419 2459 -411
rect 2500 -419 2503 -411
rect 2506 -419 2520 -411
rect 2523 -419 2527 -411
rect 572 -436 577 -429
rect 572 -440 577 -439
rect 498 -480 503 -477
rect 498 -486 503 -483
rect 572 -490 577 -487
rect 798 -487 802 -479
rect 805 -487 819 -479
rect 822 -487 825 -479
rect 954 -487 958 -479
rect 961 -487 975 -479
rect 978 -487 981 -479
rect 1104 -487 1108 -479
rect 1111 -487 1125 -479
rect 1128 -487 1131 -479
rect 1251 -487 1255 -479
rect 1258 -487 1272 -479
rect 1275 -487 1278 -479
rect 572 -496 577 -493
rect 572 -524 577 -522
rect 788 -520 796 -516
rect 838 -520 846 -516
rect 572 -534 577 -527
rect 788 -526 796 -523
rect 838 -526 846 -523
rect 944 -520 952 -516
rect 994 -520 1002 -516
rect 944 -526 952 -523
rect 994 -526 1002 -523
rect 1094 -520 1102 -516
rect 1144 -520 1152 -516
rect 1094 -526 1102 -523
rect 1144 -526 1152 -523
rect 1250 -520 1258 -516
rect 1300 -520 1308 -516
rect 1250 -526 1258 -523
rect 1300 -526 1308 -523
rect 1496 -520 1504 -516
rect 1553 -520 1561 -516
rect 1496 -526 1504 -523
rect 1553 -526 1561 -523
rect 1735 -519 1743 -515
rect 1791 -519 1799 -515
rect 1735 -525 1743 -522
rect 1791 -525 1799 -522
rect 1968 -519 1976 -515
rect 2024 -519 2032 -515
rect 1968 -525 1976 -522
rect 2024 -525 2032 -522
rect 2189 -519 2197 -515
rect 2245 -519 2253 -515
rect 2189 -525 2197 -522
rect 2245 -525 2253 -522
rect 2327 -522 2335 -518
rect 2327 -528 2335 -525
rect 572 -544 577 -537
rect 572 -548 577 -547
rect 1496 -575 1504 -572
rect 430 -586 435 -583
rect 430 -592 435 -589
rect 788 -585 796 -582
rect 572 -601 577 -598
rect 572 -607 577 -604
rect 788 -602 796 -588
rect 838 -585 846 -582
rect 944 -585 952 -582
rect 788 -609 796 -605
rect 838 -602 846 -588
rect 944 -602 952 -588
rect 994 -585 1002 -582
rect 1094 -585 1102 -582
rect 838 -609 846 -605
rect 944 -609 952 -605
rect 994 -602 1002 -588
rect 1094 -602 1102 -588
rect 1144 -585 1152 -582
rect 1250 -585 1258 -582
rect 994 -609 1002 -605
rect 1094 -609 1102 -605
rect 1144 -602 1152 -588
rect 1250 -602 1258 -588
rect 1300 -585 1308 -582
rect 1144 -609 1152 -605
rect 1250 -609 1258 -605
rect 1300 -602 1308 -588
rect 1496 -592 1504 -578
rect 1553 -575 1561 -572
rect 1735 -574 1743 -571
rect 1496 -599 1504 -595
rect 1553 -592 1561 -578
rect 1735 -591 1743 -577
rect 1791 -574 1799 -571
rect 1968 -574 1976 -571
rect 1553 -599 1561 -595
rect 1735 -598 1743 -594
rect 1791 -591 1799 -577
rect 1968 -591 1976 -577
rect 2024 -574 2032 -571
rect 2189 -574 2197 -571
rect 1791 -598 1799 -594
rect 1968 -598 1976 -594
rect 2024 -591 2032 -577
rect 2189 -591 2197 -577
rect 2245 -574 2253 -571
rect 2024 -598 2032 -594
rect 2189 -598 2197 -594
rect 2245 -591 2253 -577
rect 2327 -577 2335 -574
rect 2245 -598 2253 -594
rect 2327 -594 2335 -580
rect 2327 -601 2335 -597
rect 1300 -609 1308 -605
rect 572 -635 577 -633
rect 572 -645 577 -638
rect 572 -655 577 -648
rect 572 -659 577 -658
<< pdiffusion >>
rect 1554 304 1558 312
rect 1561 304 1575 312
rect 1578 304 1581 312
rect 1612 304 1615 312
rect 1618 304 1622 312
rect 1694 303 1695 309
rect 1698 303 1705 309
rect 1708 303 1715 309
rect 1718 303 1722 309
rect 1749 301 1752 309
rect 1755 301 1758 309
rect 1838 305 1839 311
rect 1842 305 1849 311
rect 1852 305 1859 311
rect 1862 305 1866 311
rect 1893 303 1896 311
rect 1899 303 1902 311
rect 1981 306 1982 312
rect 1985 306 1992 312
rect 1995 306 2002 312
rect 2005 306 2009 312
rect 2036 304 2039 312
rect 2042 304 2045 312
rect 968 221 969 227
rect 972 221 979 227
rect 982 221 989 227
rect 992 221 999 227
rect 1002 221 1003 227
rect 1030 219 1033 227
rect 1036 219 1039 227
rect 1099 219 1102 227
rect 1105 219 1108 227
rect 1135 221 1136 227
rect 1139 221 1146 227
rect 1149 221 1156 227
rect 1159 221 1166 227
rect 1169 221 1170 227
rect 1547 188 1550 196
rect 1553 188 1558 196
rect 1562 188 1567 196
rect 1570 188 1574 196
rect 1785 191 1788 199
rect 1791 191 1796 199
rect 1800 191 1805 199
rect 1808 191 1812 199
rect 2018 191 2021 199
rect 2024 191 2029 199
rect 2033 191 2038 199
rect 2041 191 2045 199
rect 2256 194 2259 202
rect 2262 194 2267 202
rect 2271 194 2276 202
rect 2279 194 2283 202
rect 1011 158 1019 161
rect 1339 164 1347 167
rect 1011 152 1019 155
rect 1339 158 1347 161
rect 1447 147 1455 151
rect 1142 144 1150 147
rect 1447 141 1455 144
rect 1685 150 1693 154
rect 1685 144 1693 147
rect 1918 150 1926 154
rect 1142 138 1150 141
rect 1918 144 1926 147
rect 2156 153 2164 157
rect 2156 147 2164 150
rect 2376 146 2384 150
rect 2376 140 2384 143
rect 1341 129 1346 130
rect 1013 123 1018 124
rect 798 116 806 119
rect 798 110 806 113
rect 1013 119 1018 120
rect 1341 125 1346 126
rect 1341 119 1346 120
rect 1013 113 1018 114
rect 1013 109 1018 110
rect 1144 109 1149 110
rect 1341 115 1346 116
rect 1013 103 1018 104
rect 1013 99 1018 100
rect 1144 105 1149 106
rect 1341 109 1346 110
rect 1341 105 1346 106
rect 1447 107 1455 110
rect 1532 124 1540 127
rect 1579 124 1587 127
rect 1532 116 1540 121
rect 1532 107 1540 112
rect 1579 116 1587 121
rect 1144 99 1149 100
rect 1144 95 1149 96
rect 800 81 805 82
rect 1144 89 1149 90
rect 1447 90 1455 104
rect 1532 100 1540 104
rect 1579 107 1587 112
rect 1685 110 1693 113
rect 1770 127 1778 130
rect 1817 127 1825 130
rect 1770 119 1778 124
rect 1770 110 1778 115
rect 1817 119 1825 124
rect 1579 100 1587 104
rect 1685 93 1693 107
rect 1770 103 1778 107
rect 1817 110 1825 115
rect 1817 103 1825 107
rect 1918 110 1926 113
rect 2003 127 2011 130
rect 2050 127 2058 130
rect 2003 119 2011 124
rect 2003 110 2011 115
rect 2050 119 2058 124
rect 1144 85 1149 86
rect 1447 83 1455 87
rect 1685 86 1693 90
rect 1918 93 1926 107
rect 2003 103 2011 107
rect 2050 110 2058 115
rect 2156 113 2164 116
rect 2241 130 2249 133
rect 2288 130 2296 133
rect 2450 141 2454 149
rect 2457 141 2460 149
rect 2501 141 2504 149
rect 2507 141 2512 149
rect 2516 141 2521 149
rect 2524 141 2528 149
rect 2241 122 2249 127
rect 2241 113 2249 118
rect 2288 122 2296 127
rect 2050 103 2058 107
rect 2156 96 2164 110
rect 2241 106 2249 110
rect 2288 113 2296 118
rect 2288 106 2296 110
rect 2376 96 2384 99
rect 1918 86 1926 90
rect 2156 89 2164 93
rect 2376 88 2384 93
rect 2376 79 2384 84
rect 800 77 805 78
rect 800 71 805 72
rect 800 67 805 68
rect 800 61 805 62
rect 800 57 805 58
rect 1007 62 1015 65
rect 1335 68 1343 71
rect 1007 56 1015 59
rect 1335 62 1343 65
rect 1545 60 1549 68
rect 1552 60 1557 68
rect 1561 60 1566 68
rect 1569 60 1572 68
rect 1783 63 1787 71
rect 1790 63 1795 71
rect 1799 63 1804 71
rect 1807 63 1810 71
rect 2016 63 2020 71
rect 2023 63 2028 71
rect 2032 63 2037 71
rect 2040 63 2043 71
rect 2254 66 2258 74
rect 2261 66 2266 74
rect 2270 66 2275 74
rect 2278 66 2281 74
rect 2376 72 2384 76
rect 1138 48 1146 51
rect 1138 42 1146 45
rect 794 20 802 23
rect 794 14 802 17
rect 1434 16 1442 20
rect 1434 10 1442 13
rect 1672 19 1680 23
rect 1672 13 1680 16
rect 1905 19 1913 23
rect 1905 13 1913 16
rect 2143 22 2151 26
rect 2143 16 2151 19
rect 2450 21 2454 29
rect 2457 21 2460 29
rect 2501 21 2504 29
rect 2507 21 2512 29
rect 2516 21 2521 29
rect 2524 21 2528 29
rect 854 -21 862 -18
rect 942 -16 950 -13
rect 1170 -7 1178 -4
rect 1170 -13 1178 -10
rect 1272 -9 1280 -6
rect 1272 -15 1280 -12
rect 2376 -13 2384 -9
rect 2376 -19 2384 -16
rect 854 -27 862 -24
rect 942 -22 950 -19
rect 1547 -36 1550 -28
rect 1553 -36 1558 -28
rect 1562 -36 1567 -28
rect 1570 -36 1574 -28
rect 1785 -33 1788 -25
rect 1791 -33 1796 -25
rect 1800 -33 1805 -25
rect 1808 -33 1812 -25
rect 2018 -33 2021 -25
rect 2024 -33 2029 -25
rect 2033 -33 2038 -25
rect 2041 -33 2045 -25
rect 2256 -30 2259 -22
rect 2262 -30 2267 -22
rect 2271 -30 2276 -22
rect 2279 -30 2283 -22
rect 2450 -18 2454 -10
rect 2457 -18 2460 -10
rect 2501 -18 2504 -10
rect 2507 -18 2512 -10
rect 2516 -18 2521 -10
rect 2524 -18 2528 -10
rect 1172 -42 1177 -41
rect 944 -51 949 -50
rect 856 -56 861 -55
rect 856 -60 861 -59
rect 944 -55 949 -54
rect 1172 -46 1177 -45
rect 1274 -44 1279 -43
rect 1172 -52 1177 -51
rect 944 -61 949 -60
rect 1172 -56 1177 -55
rect 1274 -48 1279 -47
rect 1434 -52 1442 -49
rect 1274 -54 1279 -53
rect 856 -66 861 -65
rect 856 -70 861 -69
rect 944 -65 949 -64
rect 856 -76 861 -75
rect 944 -71 949 -70
rect 1172 -62 1177 -61
rect 1274 -58 1279 -57
rect 1172 -66 1177 -65
rect 1274 -64 1279 -63
rect 1434 -60 1442 -55
rect 1274 -68 1279 -67
rect 1434 -69 1442 -64
rect 1672 -49 1680 -46
rect 1672 -57 1680 -52
rect 1672 -66 1680 -61
rect 1905 -49 1913 -46
rect 1905 -57 1913 -52
rect 944 -75 949 -74
rect 856 -80 861 -79
rect 1434 -76 1442 -72
rect 1672 -73 1680 -69
rect 1905 -66 1913 -61
rect 2143 -46 2151 -43
rect 2143 -54 2151 -49
rect 2143 -63 2151 -58
rect 1905 -73 1913 -69
rect 2143 -70 2151 -66
rect 2376 -63 2384 -60
rect 2376 -71 2384 -66
rect 2376 -80 2384 -75
rect 2376 -87 2384 -83
rect 850 -117 858 -114
rect 938 -112 946 -109
rect 1166 -103 1174 -100
rect 1166 -109 1174 -106
rect 1268 -105 1276 -102
rect 1268 -111 1276 -108
rect 850 -123 858 -120
rect 938 -118 946 -115
rect 1532 -100 1540 -97
rect 1579 -100 1587 -97
rect 1532 -108 1540 -103
rect 1532 -117 1540 -112
rect 1579 -108 1587 -103
rect 1435 -125 1443 -121
rect 1435 -131 1443 -128
rect 1532 -124 1540 -120
rect 1579 -117 1587 -112
rect 1770 -97 1778 -94
rect 1817 -97 1825 -94
rect 1770 -105 1778 -100
rect 1770 -114 1778 -109
rect 1817 -105 1825 -100
rect 1579 -124 1587 -120
rect 1673 -122 1681 -118
rect 1673 -128 1681 -125
rect 1770 -121 1778 -117
rect 1817 -114 1825 -109
rect 2003 -97 2011 -94
rect 2050 -97 2058 -94
rect 2003 -105 2011 -100
rect 2003 -114 2011 -109
rect 2050 -105 2058 -100
rect 1817 -121 1825 -117
rect 1906 -122 1914 -118
rect 1906 -128 1914 -125
rect 2003 -121 2011 -117
rect 2050 -114 2058 -109
rect 2241 -94 2249 -91
rect 2288 -94 2296 -91
rect 2241 -102 2249 -97
rect 2241 -111 2249 -106
rect 2288 -102 2296 -97
rect 2050 -121 2058 -117
rect 2144 -119 2152 -115
rect 2144 -125 2152 -122
rect 2241 -118 2249 -114
rect 2288 -111 2296 -106
rect 2288 -118 2296 -114
rect 2450 -138 2454 -130
rect 2457 -138 2460 -130
rect 2501 -138 2504 -130
rect 2507 -138 2512 -130
rect 2516 -138 2521 -130
rect 2524 -138 2528 -130
rect 1545 -164 1549 -156
rect 1552 -164 1557 -156
rect 1561 -164 1566 -156
rect 1569 -164 1572 -156
rect 1783 -161 1787 -153
rect 1790 -161 1795 -153
rect 1799 -161 1804 -153
rect 1807 -161 1810 -153
rect 2016 -161 2020 -153
rect 2023 -161 2028 -153
rect 2032 -161 2037 -153
rect 2040 -161 2043 -153
rect 2254 -158 2258 -150
rect 2261 -158 2266 -150
rect 2270 -158 2275 -150
rect 2278 -158 2281 -150
rect 1388 -180 1396 -176
rect 1007 -197 1015 -193
rect 1007 -203 1015 -200
rect 1157 -197 1165 -193
rect 1388 -186 1396 -183
rect 1435 -193 1443 -190
rect 1157 -203 1165 -200
rect 1304 -197 1312 -193
rect 1304 -203 1312 -200
rect 1435 -201 1443 -196
rect 1435 -210 1443 -205
rect 1673 -190 1681 -187
rect 1673 -198 1681 -193
rect 1673 -207 1681 -202
rect 1906 -190 1914 -187
rect 1906 -198 1914 -193
rect 1435 -217 1443 -213
rect 1673 -214 1681 -210
rect 1906 -207 1914 -202
rect 2144 -187 2152 -184
rect 2375 -167 2383 -163
rect 2375 -173 2383 -170
rect 2449 -172 2453 -164
rect 2456 -172 2459 -164
rect 2500 -172 2503 -164
rect 2506 -172 2511 -164
rect 2515 -172 2520 -164
rect 2523 -172 2527 -164
rect 2144 -195 2152 -190
rect 2144 -204 2152 -199
rect 1906 -214 1914 -210
rect 2144 -211 2152 -207
rect 2375 -217 2383 -214
rect 1388 -230 1396 -227
rect 2375 -225 2383 -220
rect 1007 -247 1015 -244
rect 605 -269 610 -266
rect 1007 -255 1015 -250
rect 1157 -247 1165 -244
rect 1007 -264 1015 -259
rect 605 -275 610 -272
rect 1007 -271 1015 -267
rect 1157 -255 1165 -250
rect 1304 -247 1312 -244
rect 1157 -264 1165 -259
rect 1157 -271 1165 -267
rect 1304 -255 1312 -250
rect 1388 -238 1396 -233
rect 2375 -234 2383 -229
rect 1388 -247 1396 -242
rect 2375 -241 2383 -237
rect 1388 -254 1396 -250
rect 1304 -264 1312 -259
rect 1304 -271 1312 -267
rect 1470 -268 1473 -260
rect 1476 -268 1481 -260
rect 1485 -268 1490 -260
rect 1493 -268 1497 -260
rect 1708 -265 1711 -257
rect 1714 -265 1719 -257
rect 1723 -265 1728 -257
rect 1731 -265 1735 -257
rect 1941 -265 1944 -257
rect 1947 -265 1952 -257
rect 1956 -265 1961 -257
rect 1964 -265 1968 -257
rect 2179 -262 2182 -254
rect 2185 -262 2190 -254
rect 2194 -262 2199 -254
rect 2202 -262 2206 -254
rect 792 -289 800 -285
rect 792 -295 800 -292
rect 948 -289 956 -285
rect 948 -295 956 -292
rect 1098 -289 1106 -285
rect 1098 -295 1106 -292
rect 1245 -289 1253 -285
rect 1245 -295 1253 -292
rect 2449 -292 2453 -284
rect 2456 -292 2459 -284
rect 2500 -292 2503 -284
rect 2506 -292 2511 -284
rect 2515 -292 2520 -284
rect 2523 -292 2527 -284
rect 605 -303 610 -302
rect 605 -307 610 -306
rect 605 -313 610 -312
rect 605 -317 610 -316
rect 605 -323 610 -322
rect 800 -326 803 -318
rect 806 -326 811 -318
rect 815 -326 820 -318
rect 823 -326 827 -318
rect 956 -326 959 -318
rect 962 -326 967 -318
rect 971 -326 976 -318
rect 979 -326 983 -318
rect 1106 -326 1109 -318
rect 1112 -326 1117 -318
rect 1121 -326 1126 -318
rect 1129 -326 1133 -318
rect 1253 -326 1256 -318
rect 1259 -326 1264 -318
rect 1268 -326 1273 -318
rect 1276 -326 1280 -318
rect 605 -327 610 -326
rect 667 -345 675 -341
rect 667 -362 675 -348
rect 1455 -332 1463 -329
rect 1502 -332 1510 -329
rect 1455 -340 1463 -335
rect 1455 -349 1463 -344
rect 1502 -340 1510 -335
rect 1455 -356 1463 -352
rect 1502 -349 1510 -344
rect 1693 -329 1701 -326
rect 1740 -329 1748 -326
rect 1693 -337 1701 -332
rect 1693 -346 1701 -341
rect 1740 -337 1748 -332
rect 1502 -356 1510 -352
rect 1693 -353 1701 -349
rect 1740 -346 1748 -341
rect 1926 -329 1934 -326
rect 1973 -329 1981 -326
rect 1926 -337 1934 -332
rect 1926 -346 1934 -341
rect 1973 -337 1981 -332
rect 1740 -353 1748 -349
rect 1926 -353 1934 -349
rect 1973 -346 1981 -341
rect 2164 -326 2172 -323
rect 2211 -326 2219 -323
rect 2375 -326 2383 -322
rect 2164 -334 2172 -329
rect 2164 -343 2172 -338
rect 2211 -334 2219 -329
rect 1973 -353 1981 -349
rect 2164 -350 2172 -346
rect 2211 -343 2219 -338
rect 2375 -332 2383 -329
rect 2449 -331 2453 -323
rect 2456 -331 2459 -323
rect 2500 -331 2503 -323
rect 2506 -331 2511 -323
rect 2515 -331 2520 -323
rect 2523 -331 2527 -323
rect 2211 -350 2219 -346
rect 667 -368 675 -365
rect 2375 -376 2383 -373
rect 605 -382 610 -379
rect 605 -388 610 -385
rect 667 -402 675 -399
rect 667 -409 675 -405
rect 785 -390 793 -387
rect 832 -390 840 -387
rect 785 -398 793 -393
rect 785 -407 793 -402
rect 832 -398 840 -393
rect 605 -416 610 -415
rect 785 -414 793 -410
rect 832 -407 840 -402
rect 941 -390 949 -387
rect 988 -390 996 -387
rect 941 -398 949 -393
rect 941 -407 949 -402
rect 988 -398 996 -393
rect 832 -414 840 -410
rect 941 -414 949 -410
rect 988 -407 996 -402
rect 1091 -390 1099 -387
rect 1138 -390 1146 -387
rect 1091 -398 1099 -393
rect 1091 -407 1099 -402
rect 1138 -398 1146 -393
rect 988 -414 996 -410
rect 1091 -414 1099 -410
rect 1138 -407 1146 -402
rect 1238 -390 1246 -387
rect 1285 -390 1293 -387
rect 1238 -398 1246 -393
rect 1238 -407 1246 -402
rect 1285 -398 1293 -393
rect 1138 -414 1146 -410
rect 1238 -414 1246 -410
rect 1285 -407 1293 -402
rect 1468 -396 1472 -388
rect 1475 -396 1480 -388
rect 1484 -396 1489 -388
rect 1492 -396 1495 -388
rect 1706 -393 1710 -385
rect 1713 -393 1718 -385
rect 1722 -393 1727 -385
rect 1730 -393 1733 -385
rect 1939 -393 1943 -385
rect 1946 -393 1951 -385
rect 1955 -393 1960 -385
rect 1963 -393 1966 -385
rect 2177 -390 2181 -382
rect 2184 -390 2189 -382
rect 2193 -390 2198 -382
rect 2201 -390 2204 -382
rect 2375 -384 2383 -379
rect 1285 -414 1293 -410
rect 605 -420 610 -419
rect 2375 -393 2383 -388
rect 2375 -400 2383 -396
rect 605 -426 610 -425
rect 605 -430 610 -429
rect 605 -436 610 -435
rect 605 -440 610 -439
rect 798 -454 802 -446
rect 805 -454 810 -446
rect 814 -454 819 -446
rect 822 -454 825 -446
rect 954 -454 958 -446
rect 961 -454 966 -446
rect 970 -454 975 -446
rect 978 -454 981 -446
rect 1104 -454 1108 -446
rect 1111 -454 1116 -446
rect 1120 -454 1125 -446
rect 1128 -454 1131 -446
rect 1251 -454 1255 -446
rect 1258 -454 1263 -446
rect 1267 -454 1272 -446
rect 1275 -454 1278 -446
rect 2449 -451 2453 -443
rect 2456 -451 2459 -443
rect 2500 -451 2503 -443
rect 2506 -451 2511 -443
rect 2515 -451 2520 -443
rect 2523 -451 2527 -443
rect 465 -480 470 -477
rect 465 -486 470 -483
rect 605 -490 610 -487
rect 605 -496 610 -493
rect 756 -520 764 -516
rect 605 -524 610 -523
rect 756 -526 764 -523
rect 605 -528 610 -527
rect 870 -520 878 -516
rect 912 -520 920 -516
rect 870 -526 878 -523
rect 912 -526 920 -523
rect 1026 -520 1034 -516
rect 1062 -520 1070 -516
rect 1026 -526 1034 -523
rect 1062 -526 1070 -523
rect 1176 -520 1184 -516
rect 1218 -520 1226 -516
rect 1176 -526 1184 -523
rect 1218 -526 1226 -523
rect 1332 -520 1340 -516
rect 1464 -520 1472 -516
rect 1332 -526 1340 -523
rect 1464 -526 1472 -523
rect 1585 -520 1593 -516
rect 1703 -519 1711 -515
rect 1585 -526 1593 -523
rect 1703 -525 1711 -522
rect 1823 -519 1831 -515
rect 1936 -519 1944 -515
rect 1823 -525 1831 -522
rect 1936 -525 1944 -522
rect 2056 -519 2064 -515
rect 2157 -519 2165 -515
rect 2056 -525 2064 -522
rect 2157 -525 2165 -522
rect 2277 -519 2285 -515
rect 2277 -525 2285 -522
rect 2359 -522 2367 -518
rect 2359 -528 2367 -525
rect 605 -534 610 -533
rect 605 -538 610 -537
rect 605 -544 610 -543
rect 605 -548 610 -547
rect 1464 -575 1472 -572
rect 463 -586 468 -583
rect 756 -585 764 -582
rect 463 -592 468 -589
rect 756 -593 764 -588
rect 605 -601 610 -598
rect 756 -602 764 -597
rect 870 -585 878 -582
rect 912 -585 920 -582
rect 605 -607 610 -604
rect 756 -609 764 -605
rect 870 -593 878 -588
rect 870 -602 878 -597
rect 912 -593 920 -588
rect 912 -602 920 -597
rect 1026 -585 1034 -582
rect 1062 -585 1070 -582
rect 870 -609 878 -605
rect 912 -609 920 -605
rect 1026 -593 1034 -588
rect 1026 -602 1034 -597
rect 1062 -593 1070 -588
rect 1062 -602 1070 -597
rect 1176 -585 1184 -582
rect 1218 -585 1226 -582
rect 1026 -609 1034 -605
rect 1062 -609 1070 -605
rect 1176 -593 1184 -588
rect 1176 -602 1184 -597
rect 1218 -593 1226 -588
rect 1218 -602 1226 -597
rect 1332 -585 1340 -582
rect 1464 -583 1472 -578
rect 1176 -609 1184 -605
rect 1218 -609 1226 -605
rect 1332 -593 1340 -588
rect 1464 -592 1472 -587
rect 1585 -575 1593 -572
rect 1703 -574 1711 -571
rect 1332 -602 1340 -597
rect 1464 -599 1472 -595
rect 1585 -583 1593 -578
rect 1585 -592 1593 -587
rect 1703 -582 1711 -577
rect 1703 -591 1711 -586
rect 1823 -574 1831 -571
rect 1936 -574 1944 -571
rect 1585 -599 1593 -595
rect 1703 -598 1711 -594
rect 1823 -582 1831 -577
rect 1823 -591 1831 -586
rect 1936 -582 1944 -577
rect 1936 -591 1944 -586
rect 2056 -574 2064 -571
rect 2157 -574 2165 -571
rect 1823 -598 1831 -594
rect 1936 -598 1944 -594
rect 2056 -582 2064 -577
rect 2056 -591 2064 -586
rect 2157 -582 2165 -577
rect 2157 -591 2165 -586
rect 2277 -574 2285 -571
rect 2056 -598 2064 -594
rect 2157 -598 2165 -594
rect 2277 -582 2285 -577
rect 2359 -577 2367 -574
rect 2277 -591 2285 -586
rect 2277 -598 2285 -594
rect 2359 -585 2367 -580
rect 2359 -594 2367 -589
rect 2359 -601 2367 -597
rect 1332 -609 1340 -605
rect 605 -635 610 -634
rect 605 -639 610 -638
rect 605 -645 610 -644
rect 605 -649 610 -648
rect 605 -655 610 -654
rect 605 -659 610 -658
<< ndcontact >>
rect 1550 336 1554 344
rect 1565 336 1570 344
rect 1581 336 1585 344
rect 1608 336 1612 344
rect 1622 336 1626 344
rect 1689 338 1694 344
rect 1699 338 1704 344
rect 1709 338 1714 344
rect 1719 338 1724 344
rect 1745 333 1749 341
rect 1758 333 1762 341
rect 1833 340 1838 346
rect 1843 340 1848 346
rect 1853 340 1858 346
rect 1863 340 1868 346
rect 1889 335 1893 343
rect 1902 335 1906 343
rect 1976 341 1981 347
rect 1986 341 1991 347
rect 1996 341 2001 347
rect 2006 341 2011 347
rect 2032 336 2036 344
rect 2045 336 2049 344
rect 963 256 968 262
rect 973 256 978 262
rect 983 256 988 262
rect 993 256 998 262
rect 1003 256 1008 262
rect 1026 251 1030 259
rect 1039 251 1043 259
rect 1095 251 1099 259
rect 1108 251 1112 259
rect 1130 256 1135 262
rect 1140 256 1145 262
rect 1150 256 1155 262
rect 1160 256 1165 262
rect 1170 256 1175 262
rect 1307 167 1315 171
rect 979 161 987 165
rect 979 148 987 152
rect 1307 154 1315 158
rect 1543 156 1547 164
rect 1578 156 1582 164
rect 1781 159 1785 167
rect 1816 159 1820 167
rect 2014 159 2018 167
rect 2049 159 2053 167
rect 2252 162 2256 170
rect 2287 162 2291 170
rect 1110 147 1118 151
rect 1479 151 1487 155
rect 1717 154 1725 158
rect 1950 154 1958 158
rect 1110 134 1118 138
rect 1479 137 1487 141
rect 1717 140 1725 144
rect 2188 157 2196 161
rect 1950 140 1958 144
rect 2188 143 2196 147
rect 2408 150 2416 154
rect 1308 130 1313 135
rect 980 124 985 129
rect 766 119 774 123
rect 1500 127 1508 131
rect 766 106 774 110
rect 1111 110 1116 115
rect 980 94 985 99
rect 1308 100 1313 105
rect 1479 110 1487 114
rect 1611 127 1619 131
rect 1738 130 1746 134
rect 767 82 772 87
rect 1479 94 1487 99
rect 1500 96 1508 100
rect 1717 113 1725 117
rect 1849 130 1857 134
rect 1971 130 1979 134
rect 1611 96 1619 100
rect 1717 97 1725 102
rect 1738 99 1746 103
rect 1950 113 1958 117
rect 2082 130 2090 134
rect 2209 133 2217 137
rect 1849 99 1857 103
rect 1111 80 1116 85
rect 1479 79 1487 83
rect 1950 97 1958 102
rect 1971 99 1979 103
rect 2188 116 2196 120
rect 2320 133 2328 137
rect 2408 136 2416 140
rect 2082 99 2090 103
rect 2188 100 2196 105
rect 2209 102 2217 106
rect 2446 109 2450 117
rect 2460 109 2464 117
rect 2497 109 2501 117
rect 2528 109 2532 117
rect 2320 102 2328 106
rect 2408 99 2416 103
rect 1717 82 1725 86
rect 1950 82 1958 86
rect 2188 85 2196 89
rect 1303 71 1311 75
rect 975 65 983 69
rect 767 52 772 57
rect 975 52 983 56
rect 1303 58 1311 62
rect 2408 68 2416 72
rect 1106 51 1114 55
rect 1106 38 1114 42
rect 2446 53 2450 61
rect 2460 53 2464 61
rect 2497 53 2501 61
rect 2528 53 2532 61
rect 1541 27 1545 35
rect 1572 27 1576 35
rect 1779 30 1783 38
rect 1810 30 1814 38
rect 2012 30 2016 38
rect 2043 30 2047 38
rect 2250 33 2254 41
rect 2281 33 2285 41
rect 762 23 770 27
rect 762 10 770 14
rect 1466 20 1474 24
rect 1704 23 1712 27
rect 1937 23 1945 27
rect 1466 6 1474 10
rect 1704 9 1712 13
rect 2175 26 2183 30
rect 1937 9 1945 13
rect 2175 12 2183 16
rect 1138 -4 1146 0
rect 910 -13 918 -9
rect 822 -18 830 -14
rect 1240 -6 1248 -2
rect 1138 -17 1146 -13
rect 1240 -19 1248 -15
rect 2408 -9 2416 -5
rect 822 -31 830 -27
rect 910 -26 918 -22
rect 2408 -23 2416 -19
rect 1139 -41 1144 -36
rect 911 -50 916 -45
rect 1241 -43 1246 -38
rect 823 -55 828 -50
rect 1466 -49 1474 -45
rect 1139 -71 1144 -66
rect 1241 -73 1246 -68
rect 1704 -46 1712 -42
rect 1543 -68 1547 -60
rect 1578 -68 1582 -60
rect 1937 -46 1945 -42
rect 1781 -65 1785 -57
rect 1816 -65 1820 -57
rect 911 -80 916 -75
rect 1466 -80 1474 -76
rect 2175 -43 2183 -39
rect 2014 -65 2018 -57
rect 2049 -65 2053 -57
rect 2446 -50 2450 -42
rect 2460 -50 2464 -42
rect 2497 -50 2501 -42
rect 2528 -50 2532 -42
rect 2252 -62 2256 -54
rect 2287 -62 2291 -54
rect 1704 -77 1712 -73
rect 1937 -77 1945 -73
rect 2408 -60 2416 -56
rect 2175 -74 2183 -70
rect 823 -85 828 -80
rect 1134 -100 1142 -96
rect 1500 -97 1508 -93
rect 906 -109 914 -105
rect 818 -114 826 -110
rect 1236 -102 1244 -98
rect 1134 -113 1142 -109
rect 1236 -115 1244 -111
rect 818 -127 826 -123
rect 906 -122 914 -118
rect 1611 -97 1619 -93
rect 1738 -94 1746 -90
rect 1467 -121 1475 -117
rect 1500 -128 1508 -124
rect 1849 -94 1857 -90
rect 1971 -94 1979 -90
rect 1705 -118 1713 -114
rect 1611 -128 1619 -124
rect 1738 -125 1746 -121
rect 2082 -94 2090 -90
rect 2209 -91 2217 -87
rect 1849 -125 1857 -121
rect 1938 -118 1946 -114
rect 1467 -135 1475 -131
rect 1705 -132 1713 -128
rect 1971 -125 1979 -121
rect 2320 -91 2328 -87
rect 2408 -91 2416 -87
rect 2176 -115 2184 -111
rect 2082 -125 2090 -121
rect 2209 -122 2217 -118
rect 2446 -106 2450 -98
rect 2460 -106 2464 -98
rect 2497 -106 2501 -98
rect 2528 -106 2532 -98
rect 2320 -122 2328 -118
rect 1938 -132 1946 -128
rect 2176 -129 2184 -125
rect 1356 -176 1364 -172
rect 975 -193 983 -189
rect 1125 -193 1133 -189
rect 975 -207 983 -203
rect 1272 -193 1280 -189
rect 1356 -190 1364 -186
rect 1467 -190 1475 -186
rect 1125 -207 1133 -203
rect 1272 -207 1280 -203
rect 1541 -197 1545 -189
rect 1572 -197 1576 -189
rect 1705 -187 1713 -183
rect 1779 -194 1783 -186
rect 1810 -194 1814 -186
rect 1938 -187 1946 -183
rect 1467 -221 1475 -217
rect 2012 -194 2016 -186
rect 2043 -194 2047 -186
rect 2176 -184 2184 -180
rect 2407 -163 2415 -159
rect 2407 -177 2415 -173
rect 2250 -191 2254 -183
rect 2281 -191 2285 -183
rect 1705 -218 1713 -214
rect 1938 -218 1946 -214
rect 2445 -204 2449 -196
rect 2459 -204 2463 -196
rect 2496 -204 2500 -196
rect 2527 -204 2531 -196
rect 2176 -215 2184 -211
rect 2407 -214 2415 -210
rect 1356 -227 1364 -223
rect 975 -244 983 -240
rect 1125 -244 1133 -240
rect 572 -266 577 -262
rect 1272 -244 1280 -240
rect 572 -279 577 -275
rect 975 -275 983 -271
rect 1125 -275 1133 -271
rect 2407 -245 2415 -241
rect 1356 -258 1364 -254
rect 1272 -275 1280 -271
rect 2445 -260 2449 -252
rect 2459 -260 2463 -252
rect 2496 -260 2500 -252
rect 2527 -260 2531 -252
rect 760 -285 768 -281
rect 916 -285 924 -281
rect 572 -301 577 -297
rect 760 -299 768 -295
rect 1066 -285 1074 -281
rect 916 -299 924 -295
rect 1213 -285 1221 -281
rect 1066 -299 1074 -295
rect 1213 -299 1221 -295
rect 1466 -300 1470 -292
rect 1501 -300 1505 -292
rect 1704 -297 1708 -289
rect 1739 -297 1743 -289
rect 1937 -297 1941 -289
rect 1972 -297 1976 -289
rect 2175 -294 2179 -286
rect 2210 -294 2214 -286
rect 572 -332 577 -327
rect 699 -341 707 -337
rect 1423 -329 1431 -325
rect 1534 -329 1542 -325
rect 1661 -326 1669 -322
rect 699 -357 707 -352
rect 796 -358 800 -350
rect 831 -358 835 -350
rect 952 -358 956 -350
rect 987 -358 991 -350
rect 1102 -358 1106 -350
rect 1137 -358 1141 -350
rect 1249 -358 1253 -350
rect 1284 -358 1288 -350
rect 1423 -360 1431 -356
rect 1772 -326 1780 -322
rect 1894 -326 1902 -322
rect 1534 -360 1542 -356
rect 1661 -357 1669 -353
rect 2005 -326 2013 -322
rect 2132 -323 2140 -319
rect 1772 -357 1780 -353
rect 1894 -357 1902 -353
rect 2243 -323 2251 -319
rect 2407 -322 2415 -318
rect 2005 -357 2013 -353
rect 2132 -354 2140 -350
rect 2407 -336 2415 -332
rect 2243 -354 2251 -350
rect 2445 -363 2449 -355
rect 2459 -363 2463 -355
rect 2496 -363 2500 -355
rect 2527 -363 2531 -355
rect 699 -372 707 -368
rect 572 -379 577 -375
rect 2407 -373 2415 -369
rect 572 -392 577 -388
rect 753 -387 761 -383
rect 699 -399 707 -395
rect 572 -414 577 -410
rect 864 -387 872 -383
rect 909 -387 917 -383
rect 699 -413 707 -409
rect 753 -418 761 -414
rect 1020 -387 1028 -383
rect 1059 -387 1067 -383
rect 864 -418 872 -414
rect 909 -418 917 -414
rect 1170 -387 1178 -383
rect 1206 -387 1214 -383
rect 1020 -418 1028 -414
rect 1059 -418 1067 -414
rect 1317 -387 1325 -383
rect 1170 -418 1178 -414
rect 1206 -418 1214 -414
rect 1317 -418 1325 -414
rect 2407 -404 2415 -400
rect 1464 -429 1468 -421
rect 1495 -429 1499 -421
rect 1702 -426 1706 -418
rect 1733 -426 1737 -418
rect 1935 -426 1939 -418
rect 1966 -426 1970 -418
rect 2173 -423 2177 -415
rect 2204 -423 2208 -415
rect 2445 -419 2449 -411
rect 2459 -419 2463 -411
rect 2496 -419 2500 -411
rect 2527 -419 2531 -411
rect 572 -445 577 -440
rect 498 -477 503 -473
rect 498 -490 503 -486
rect 572 -487 577 -483
rect 794 -487 798 -479
rect 825 -487 829 -479
rect 950 -487 954 -479
rect 981 -487 985 -479
rect 1100 -487 1104 -479
rect 1131 -487 1135 -479
rect 1247 -487 1251 -479
rect 1278 -487 1282 -479
rect 572 -500 577 -496
rect 572 -522 577 -518
rect 788 -516 796 -512
rect 838 -516 846 -512
rect 788 -530 796 -526
rect 944 -516 952 -512
rect 838 -530 846 -526
rect 994 -516 1002 -512
rect 944 -530 952 -526
rect 1094 -516 1102 -512
rect 994 -530 1002 -526
rect 1144 -516 1152 -512
rect 1094 -530 1102 -526
rect 1250 -516 1258 -512
rect 1144 -530 1152 -526
rect 1300 -516 1308 -512
rect 1250 -530 1258 -526
rect 1496 -516 1504 -512
rect 1300 -530 1308 -526
rect 1553 -516 1561 -512
rect 1496 -530 1504 -526
rect 1735 -515 1743 -511
rect 1553 -530 1561 -526
rect 1791 -515 1799 -511
rect 1735 -529 1743 -525
rect 1968 -515 1976 -511
rect 1791 -529 1799 -525
rect 2024 -515 2032 -511
rect 1968 -529 1976 -525
rect 2189 -515 2197 -511
rect 2024 -529 2032 -525
rect 2245 -515 2253 -511
rect 2189 -529 2197 -525
rect 2327 -518 2335 -514
rect 2245 -529 2253 -525
rect 2327 -532 2335 -528
rect 572 -553 577 -548
rect 1496 -572 1504 -568
rect 1553 -572 1561 -568
rect 430 -583 435 -579
rect 788 -582 796 -578
rect 838 -582 846 -578
rect 430 -596 435 -592
rect 572 -598 577 -594
rect 944 -582 952 -578
rect 994 -582 1002 -578
rect 572 -611 577 -607
rect 1094 -582 1102 -578
rect 1144 -582 1152 -578
rect 788 -613 796 -609
rect 838 -613 846 -609
rect 1250 -582 1258 -578
rect 1300 -582 1308 -578
rect 944 -613 952 -609
rect 994 -613 1002 -609
rect 1094 -613 1102 -609
rect 1144 -613 1152 -609
rect 1735 -571 1743 -567
rect 1791 -571 1799 -567
rect 1968 -571 1976 -567
rect 2024 -571 2032 -567
rect 1496 -603 1504 -599
rect 1553 -603 1561 -599
rect 2189 -571 2197 -567
rect 2245 -571 2253 -567
rect 1735 -602 1743 -598
rect 1791 -602 1799 -598
rect 2327 -574 2335 -570
rect 1968 -602 1976 -598
rect 2024 -602 2032 -598
rect 2189 -602 2197 -598
rect 2245 -602 2253 -598
rect 2327 -605 2335 -601
rect 1250 -613 1258 -609
rect 1300 -613 1308 -609
rect 572 -633 577 -629
rect 572 -664 577 -659
<< pdcontact >>
rect 1550 304 1554 312
rect 1581 304 1585 312
rect 1608 304 1612 312
rect 1622 304 1626 312
rect 1689 303 1694 309
rect 1722 303 1727 309
rect 1745 301 1749 309
rect 1758 301 1762 309
rect 1833 305 1838 311
rect 1866 305 1871 311
rect 1889 303 1893 311
rect 1902 303 1906 311
rect 1976 306 1981 312
rect 2009 306 2014 312
rect 2032 304 2036 312
rect 2045 304 2049 312
rect 963 221 968 227
rect 1003 221 1008 227
rect 1026 219 1030 227
rect 1039 219 1043 227
rect 1095 219 1099 227
rect 1108 219 1112 227
rect 1130 221 1135 227
rect 1170 221 1175 227
rect 1543 188 1547 196
rect 1558 188 1562 196
rect 1574 188 1578 196
rect 1781 191 1785 199
rect 1796 191 1800 199
rect 1812 191 1816 199
rect 2014 191 2018 199
rect 2029 191 2033 199
rect 2045 191 2049 199
rect 2252 194 2256 202
rect 2267 194 2271 202
rect 2283 194 2287 202
rect 1011 161 1019 165
rect 1339 167 1347 171
rect 1339 154 1347 158
rect 1011 148 1019 152
rect 1447 151 1455 155
rect 1142 147 1150 151
rect 1685 154 1693 158
rect 1918 154 1926 158
rect 2156 157 2164 161
rect 1142 134 1150 138
rect 1447 137 1455 141
rect 1685 140 1693 144
rect 2376 150 2384 154
rect 1918 140 1926 144
rect 2156 143 2164 147
rect 798 119 806 123
rect 1013 124 1018 128
rect 1341 130 1346 134
rect 798 106 806 110
rect 1013 114 1018 119
rect 1341 120 1346 125
rect 1532 127 1540 131
rect 1013 104 1018 109
rect 1144 110 1149 114
rect 1341 110 1346 115
rect 1013 94 1018 99
rect 1144 100 1149 105
rect 1447 110 1455 114
rect 1341 100 1346 105
rect 1579 127 1587 131
rect 1770 130 1778 134
rect 1532 112 1540 116
rect 1579 112 1587 116
rect 1144 90 1149 95
rect 800 82 805 86
rect 1685 113 1693 117
rect 1817 130 1825 134
rect 2003 130 2011 134
rect 1770 115 1778 119
rect 1817 115 1825 119
rect 1532 96 1540 100
rect 1579 96 1587 100
rect 1918 113 1926 117
rect 1770 99 1778 103
rect 1817 99 1825 103
rect 2050 130 2058 134
rect 2241 133 2249 137
rect 2003 115 2011 119
rect 2050 115 2058 119
rect 1144 80 1149 85
rect 1447 79 1455 83
rect 1685 82 1693 86
rect 2156 116 2164 120
rect 2288 133 2296 137
rect 2376 136 2384 140
rect 2446 141 2450 149
rect 2460 141 2464 149
rect 2497 141 2501 149
rect 2512 141 2516 149
rect 2528 141 2532 149
rect 2241 118 2249 122
rect 2288 118 2296 122
rect 2003 99 2011 103
rect 2050 99 2058 103
rect 2241 102 2249 106
rect 2288 102 2296 106
rect 2376 99 2384 103
rect 1918 82 1926 86
rect 2156 85 2164 89
rect 2376 84 2384 88
rect 800 72 805 77
rect 800 62 805 67
rect 1007 65 1015 69
rect 1335 71 1343 75
rect 800 52 805 57
rect 1335 58 1343 62
rect 1541 60 1545 68
rect 1557 60 1561 68
rect 1572 60 1576 68
rect 1779 63 1783 71
rect 1795 63 1799 71
rect 1810 63 1814 71
rect 2012 63 2016 71
rect 2028 63 2032 71
rect 2043 63 2047 71
rect 2250 66 2254 74
rect 2266 66 2270 74
rect 2281 66 2285 74
rect 2376 68 2384 72
rect 1007 52 1015 56
rect 1138 51 1146 55
rect 1138 38 1146 42
rect 794 23 802 27
rect 1434 20 1442 24
rect 1672 23 1680 27
rect 794 10 802 14
rect 1905 23 1913 27
rect 2143 26 2151 30
rect 1434 6 1442 10
rect 1672 9 1680 13
rect 2446 21 2450 29
rect 2460 21 2464 29
rect 2497 21 2501 29
rect 2512 21 2516 29
rect 2528 21 2532 29
rect 1905 9 1913 13
rect 2143 12 2151 16
rect 1170 -4 1178 0
rect 854 -18 862 -14
rect 942 -13 950 -9
rect 1272 -6 1280 -2
rect 1170 -17 1178 -13
rect 2376 -9 2384 -5
rect 1272 -19 1280 -15
rect 942 -26 950 -22
rect 854 -31 862 -27
rect 1543 -36 1547 -28
rect 1558 -36 1562 -28
rect 1574 -36 1578 -28
rect 1781 -33 1785 -25
rect 1796 -33 1800 -25
rect 1812 -33 1816 -25
rect 2014 -33 2018 -25
rect 2029 -33 2033 -25
rect 2045 -33 2049 -25
rect 2252 -30 2256 -22
rect 2267 -30 2271 -22
rect 2283 -30 2287 -22
rect 2376 -23 2384 -19
rect 2446 -18 2450 -10
rect 2460 -18 2464 -10
rect 2497 -18 2501 -10
rect 2512 -18 2516 -10
rect 2528 -18 2532 -10
rect 1172 -41 1177 -37
rect 856 -55 861 -51
rect 944 -50 949 -46
rect 856 -65 861 -60
rect 944 -60 949 -55
rect 1172 -51 1177 -46
rect 1274 -43 1279 -39
rect 1172 -61 1177 -56
rect 1274 -53 1279 -48
rect 1434 -49 1442 -45
rect 856 -75 861 -70
rect 944 -70 949 -65
rect 1274 -63 1279 -58
rect 1172 -71 1177 -66
rect 1434 -64 1442 -60
rect 1274 -73 1279 -68
rect 1672 -46 1680 -42
rect 1672 -61 1680 -57
rect 1905 -46 1913 -42
rect 1905 -61 1913 -57
rect 944 -80 949 -75
rect 1434 -80 1442 -76
rect 1672 -77 1680 -73
rect 2143 -43 2151 -39
rect 2143 -58 2151 -54
rect 2376 -60 2384 -56
rect 1905 -77 1913 -73
rect 2143 -74 2151 -70
rect 2376 -75 2384 -71
rect 856 -85 861 -80
rect 1166 -100 1174 -96
rect 850 -114 858 -110
rect 938 -109 946 -105
rect 1268 -102 1276 -98
rect 1532 -97 1540 -93
rect 1166 -113 1174 -109
rect 1268 -115 1276 -111
rect 1579 -97 1587 -93
rect 1770 -94 1778 -90
rect 1532 -112 1540 -108
rect 1579 -112 1587 -108
rect 938 -122 946 -118
rect 1435 -121 1443 -117
rect 850 -127 858 -123
rect 1817 -94 1825 -90
rect 2003 -94 2011 -90
rect 1770 -109 1778 -105
rect 1817 -109 1825 -105
rect 1673 -118 1681 -114
rect 1532 -128 1540 -124
rect 1579 -128 1587 -124
rect 2050 -94 2058 -90
rect 2241 -91 2249 -87
rect 2003 -109 2011 -105
rect 2050 -109 2058 -105
rect 1770 -125 1778 -121
rect 1817 -125 1825 -121
rect 1906 -118 1914 -114
rect 1435 -135 1443 -131
rect 1673 -132 1681 -128
rect 2288 -91 2296 -87
rect 2376 -91 2384 -87
rect 2241 -106 2249 -102
rect 2288 -106 2296 -102
rect 2144 -115 2152 -111
rect 2003 -125 2011 -121
rect 2050 -125 2058 -121
rect 2241 -122 2249 -118
rect 2288 -122 2296 -118
rect 1906 -132 1914 -128
rect 2144 -129 2152 -125
rect 2446 -138 2450 -130
rect 2460 -138 2464 -130
rect 2497 -138 2501 -130
rect 2512 -138 2516 -130
rect 2528 -138 2532 -130
rect 1541 -164 1545 -156
rect 1557 -164 1561 -156
rect 1572 -164 1576 -156
rect 1779 -161 1783 -153
rect 1795 -161 1799 -153
rect 1810 -161 1814 -153
rect 2012 -161 2016 -153
rect 2028 -161 2032 -153
rect 2043 -161 2047 -153
rect 2250 -158 2254 -150
rect 2266 -158 2270 -150
rect 2281 -158 2285 -150
rect 1388 -176 1396 -172
rect 1007 -193 1015 -189
rect 1157 -193 1165 -189
rect 1007 -207 1015 -203
rect 1304 -193 1312 -189
rect 1388 -190 1396 -186
rect 1435 -190 1443 -186
rect 1673 -187 1681 -183
rect 1157 -207 1165 -203
rect 1304 -207 1312 -203
rect 1435 -205 1443 -201
rect 1673 -202 1681 -198
rect 1906 -187 1914 -183
rect 2144 -184 2152 -180
rect 1906 -202 1914 -198
rect 1435 -221 1443 -217
rect 1673 -218 1681 -214
rect 2375 -163 2383 -159
rect 2375 -177 2383 -173
rect 2445 -172 2449 -164
rect 2459 -172 2463 -164
rect 2496 -172 2500 -164
rect 2511 -172 2515 -164
rect 2527 -172 2531 -164
rect 2144 -199 2152 -195
rect 1906 -218 1914 -214
rect 2144 -215 2152 -211
rect 2375 -214 2383 -210
rect 1388 -227 1396 -223
rect 2375 -229 2383 -225
rect 1007 -244 1015 -240
rect 605 -266 610 -262
rect 1157 -244 1165 -240
rect 1007 -259 1015 -255
rect 1304 -244 1312 -240
rect 1157 -259 1165 -255
rect 1007 -275 1015 -271
rect 1388 -242 1396 -238
rect 2375 -245 2383 -241
rect 1304 -259 1312 -255
rect 1388 -258 1396 -254
rect 1157 -275 1165 -271
rect 1466 -268 1470 -260
rect 1481 -268 1485 -260
rect 1497 -268 1501 -260
rect 1704 -265 1708 -257
rect 1719 -265 1723 -257
rect 1735 -265 1739 -257
rect 1937 -265 1941 -257
rect 1952 -265 1956 -257
rect 1968 -265 1972 -257
rect 2175 -262 2179 -254
rect 2190 -262 2194 -254
rect 2206 -262 2210 -254
rect 1304 -275 1312 -271
rect 605 -279 610 -275
rect 792 -285 800 -281
rect 948 -285 956 -281
rect 605 -302 610 -298
rect 792 -299 800 -295
rect 1098 -285 1106 -281
rect 948 -299 956 -295
rect 1245 -285 1253 -281
rect 1098 -299 1106 -295
rect 1245 -299 1253 -295
rect 2445 -292 2449 -284
rect 2459 -292 2463 -284
rect 2496 -292 2500 -284
rect 2511 -292 2515 -284
rect 2527 -292 2531 -284
rect 605 -312 610 -307
rect 605 -322 610 -317
rect 796 -326 800 -318
rect 811 -326 815 -318
rect 827 -326 831 -318
rect 952 -326 956 -318
rect 967 -326 971 -318
rect 983 -326 987 -318
rect 1102 -326 1106 -318
rect 1117 -326 1121 -318
rect 1133 -326 1137 -318
rect 1249 -326 1253 -318
rect 1264 -326 1268 -318
rect 1280 -326 1284 -318
rect 605 -332 610 -327
rect 667 -341 675 -337
rect 1455 -329 1463 -325
rect 1502 -329 1510 -325
rect 1693 -326 1701 -322
rect 1455 -344 1463 -340
rect 1502 -344 1510 -340
rect 1740 -326 1748 -322
rect 1926 -326 1934 -322
rect 1693 -341 1701 -337
rect 1740 -341 1748 -337
rect 1455 -360 1463 -356
rect 1502 -360 1510 -356
rect 1973 -326 1981 -322
rect 2164 -323 2172 -319
rect 1926 -341 1934 -337
rect 1973 -341 1981 -337
rect 1693 -357 1701 -353
rect 1740 -357 1748 -353
rect 2211 -323 2219 -319
rect 2375 -322 2383 -318
rect 2164 -338 2172 -334
rect 2211 -338 2219 -334
rect 1926 -357 1934 -353
rect 1973 -357 1981 -353
rect 2375 -336 2383 -332
rect 2445 -331 2449 -323
rect 2459 -331 2463 -323
rect 2496 -331 2500 -323
rect 2511 -331 2515 -323
rect 2527 -331 2531 -323
rect 2164 -354 2172 -350
rect 2211 -354 2219 -350
rect 667 -372 675 -368
rect 2375 -373 2383 -369
rect 605 -379 610 -375
rect 605 -392 610 -388
rect 785 -387 793 -383
rect 667 -399 675 -395
rect 605 -415 610 -411
rect 667 -413 675 -409
rect 832 -387 840 -383
rect 941 -387 949 -383
rect 785 -402 793 -398
rect 832 -402 840 -398
rect 988 -387 996 -383
rect 1091 -387 1099 -383
rect 941 -402 949 -398
rect 988 -402 996 -398
rect 785 -418 793 -414
rect 832 -418 840 -414
rect 1138 -387 1146 -383
rect 1238 -387 1246 -383
rect 1091 -402 1099 -398
rect 1138 -402 1146 -398
rect 941 -418 949 -414
rect 988 -418 996 -414
rect 1285 -387 1293 -383
rect 1238 -402 1246 -398
rect 1285 -402 1293 -398
rect 1091 -418 1099 -414
rect 1138 -418 1146 -414
rect 1464 -396 1468 -388
rect 1480 -396 1484 -388
rect 1495 -396 1499 -388
rect 1702 -393 1706 -385
rect 1718 -393 1722 -385
rect 1733 -393 1737 -385
rect 1935 -393 1939 -385
rect 1951 -393 1955 -385
rect 1966 -393 1970 -385
rect 2173 -390 2177 -382
rect 2189 -390 2193 -382
rect 2204 -390 2208 -382
rect 2375 -388 2383 -384
rect 1238 -418 1246 -414
rect 1285 -418 1293 -414
rect 605 -425 610 -420
rect 2375 -404 2383 -400
rect 605 -435 610 -430
rect 605 -445 610 -440
rect 794 -454 798 -446
rect 810 -454 814 -446
rect 825 -454 829 -446
rect 950 -454 954 -446
rect 966 -454 970 -446
rect 981 -454 985 -446
rect 1100 -454 1104 -446
rect 1116 -454 1120 -446
rect 1131 -454 1135 -446
rect 1247 -454 1251 -446
rect 1263 -454 1267 -446
rect 1278 -454 1282 -446
rect 2445 -451 2449 -443
rect 2459 -451 2463 -443
rect 2496 -451 2500 -443
rect 2511 -451 2515 -443
rect 2527 -451 2531 -443
rect 465 -477 470 -473
rect 465 -490 470 -486
rect 605 -487 610 -483
rect 605 -500 610 -496
rect 756 -516 764 -512
rect 605 -523 610 -519
rect 870 -516 878 -512
rect 605 -533 610 -528
rect 756 -530 764 -526
rect 912 -516 920 -512
rect 870 -530 878 -526
rect 1026 -516 1034 -512
rect 912 -530 920 -526
rect 1062 -516 1070 -512
rect 1026 -530 1034 -526
rect 1176 -516 1184 -512
rect 1062 -530 1070 -526
rect 1218 -516 1226 -512
rect 1176 -530 1184 -526
rect 1332 -516 1340 -512
rect 1218 -530 1226 -526
rect 1464 -516 1472 -512
rect 1332 -530 1340 -526
rect 1585 -516 1593 -512
rect 1464 -530 1472 -526
rect 1703 -515 1711 -511
rect 1585 -530 1593 -526
rect 1823 -515 1831 -511
rect 1703 -529 1711 -525
rect 1936 -515 1944 -511
rect 1823 -529 1831 -525
rect 2056 -515 2064 -511
rect 1936 -529 1944 -525
rect 2157 -515 2165 -511
rect 2056 -529 2064 -525
rect 2277 -515 2285 -511
rect 2157 -529 2165 -525
rect 2359 -518 2367 -514
rect 2277 -529 2285 -525
rect 2359 -532 2367 -528
rect 605 -543 610 -538
rect 605 -553 610 -548
rect 1464 -572 1472 -568
rect 463 -583 468 -579
rect 756 -582 764 -578
rect 463 -596 468 -592
rect 605 -598 610 -594
rect 756 -597 764 -593
rect 870 -582 878 -578
rect 912 -582 920 -578
rect 605 -611 610 -607
rect 756 -613 764 -609
rect 870 -597 878 -593
rect 912 -597 920 -593
rect 1026 -582 1034 -578
rect 1062 -582 1070 -578
rect 870 -613 878 -609
rect 912 -613 920 -609
rect 1026 -597 1034 -593
rect 1062 -597 1070 -593
rect 1176 -582 1184 -578
rect 1218 -582 1226 -578
rect 1026 -613 1034 -609
rect 1062 -613 1070 -609
rect 1176 -597 1184 -593
rect 1218 -597 1226 -593
rect 1332 -582 1340 -578
rect 1464 -587 1472 -583
rect 1176 -613 1184 -609
rect 1218 -613 1226 -609
rect 1585 -572 1593 -568
rect 1703 -571 1711 -567
rect 1332 -597 1340 -593
rect 1464 -603 1472 -599
rect 1585 -587 1593 -583
rect 1703 -586 1711 -582
rect 1823 -571 1831 -567
rect 1936 -571 1944 -567
rect 1585 -603 1593 -599
rect 1703 -602 1711 -598
rect 1823 -586 1831 -582
rect 1936 -586 1944 -582
rect 2056 -571 2064 -567
rect 2157 -571 2165 -567
rect 1823 -602 1831 -598
rect 1936 -602 1944 -598
rect 2056 -586 2064 -582
rect 2157 -586 2165 -582
rect 2277 -571 2285 -567
rect 2056 -602 2064 -598
rect 2157 -602 2165 -598
rect 2359 -574 2367 -570
rect 2277 -586 2285 -582
rect 2359 -589 2367 -585
rect 2277 -602 2285 -598
rect 2359 -605 2367 -601
rect 1332 -613 1340 -609
rect 605 -634 610 -630
rect 605 -644 610 -639
rect 605 -654 610 -649
rect 605 -664 610 -659
<< polysilicon >>
rect 1558 344 1561 347
rect 1575 344 1578 347
rect 1615 344 1618 347
rect 1695 344 1698 347
rect 1705 344 1708 347
rect 1715 344 1718 347
rect 1839 346 1842 349
rect 1849 346 1852 349
rect 1859 346 1862 349
rect 1982 347 1985 350
rect 1992 347 1995 350
rect 2002 347 2005 350
rect 1752 341 1755 344
rect 1558 312 1561 336
rect 1575 312 1578 336
rect 1615 332 1618 336
rect 1615 312 1618 327
rect 1695 309 1698 338
rect 1705 309 1708 338
rect 1715 309 1718 338
rect 1896 343 1899 346
rect 1752 327 1755 333
rect 1752 309 1755 322
rect 1839 311 1842 340
rect 1849 311 1852 340
rect 1859 311 1862 340
rect 2039 344 2042 347
rect 1896 329 1899 335
rect 1896 311 1899 324
rect 1982 312 1985 341
rect 1992 312 1995 341
rect 2002 312 2005 341
rect 2039 330 2042 336
rect 2039 312 2042 325
rect 1558 291 1561 304
rect 1575 291 1578 304
rect 1615 301 1618 304
rect 1695 296 1698 303
rect 1705 296 1708 303
rect 1715 296 1718 303
rect 1752 298 1755 301
rect 1839 298 1842 305
rect 1849 298 1852 305
rect 1859 298 1862 305
rect 1896 300 1899 303
rect 1982 299 1985 306
rect 1992 299 1995 306
rect 2002 299 2005 306
rect 2039 301 2042 304
rect 969 262 972 265
rect 979 262 982 265
rect 989 262 992 265
rect 999 262 1002 265
rect 1136 262 1139 265
rect 1146 262 1149 265
rect 1156 262 1159 265
rect 1166 262 1169 265
rect 1033 259 1036 262
rect 1102 259 1105 262
rect 969 227 972 256
rect 979 227 982 256
rect 989 227 992 256
rect 999 227 1002 256
rect 1033 245 1036 251
rect 1102 245 1105 251
rect 1033 227 1036 240
rect 1102 227 1105 240
rect 1136 227 1139 256
rect 1146 227 1149 256
rect 1156 227 1159 256
rect 1166 227 1169 256
rect 969 214 972 221
rect 979 214 982 221
rect 989 214 992 221
rect 999 214 1002 221
rect 1033 216 1036 219
rect 1102 216 1105 219
rect 1136 214 1139 221
rect 1146 214 1149 221
rect 1156 214 1159 221
rect 1166 214 1169 221
rect 2259 202 2262 205
rect 2276 202 2279 205
rect 1788 199 1791 202
rect 1805 199 1808 202
rect 2021 199 2024 202
rect 2038 199 2041 202
rect 1550 196 1553 199
rect 1567 196 1570 199
rect 1304 161 1307 164
rect 1315 161 1321 164
rect 976 155 979 158
rect 987 155 993 158
rect 1550 164 1553 188
rect 1567 164 1570 188
rect 1788 167 1791 191
rect 1805 167 1808 191
rect 2021 167 2024 191
rect 2038 167 2041 191
rect 2259 170 2262 194
rect 2276 170 2279 194
rect 1326 161 1339 164
rect 1347 161 1350 164
rect 998 155 1011 158
rect 1019 155 1022 158
rect 1550 153 1553 156
rect 1567 153 1570 156
rect 1107 141 1110 144
rect 1118 141 1124 144
rect 1444 144 1447 147
rect 1455 144 1470 147
rect 1129 141 1142 144
rect 1150 141 1153 144
rect 1788 156 1791 159
rect 1805 156 1808 159
rect 1682 147 1685 150
rect 1693 147 1708 150
rect 1475 144 1479 147
rect 1487 144 1490 147
rect 2021 156 2024 159
rect 2038 156 2041 159
rect 1713 147 1717 150
rect 1725 147 1728 150
rect 1915 147 1918 150
rect 1926 147 1941 150
rect 2259 159 2262 162
rect 2276 159 2279 162
rect 2153 150 2156 153
rect 2164 150 2179 153
rect 1946 147 1950 150
rect 1958 147 1961 150
rect 2184 150 2188 153
rect 2196 150 2199 153
rect 2373 143 2376 146
rect 2384 143 2399 146
rect 2454 149 2457 152
rect 2504 149 2507 152
rect 2521 149 2524 152
rect 2404 143 2408 146
rect 2416 143 2419 146
rect 1305 126 1308 129
rect 1313 126 1341 129
rect 1346 126 1349 129
rect 977 120 980 123
rect 985 120 1013 123
rect 1018 120 1021 123
rect 763 113 766 116
rect 774 113 780 116
rect 785 113 798 116
rect 806 113 809 116
rect 1497 121 1500 124
rect 1508 121 1511 124
rect 1305 116 1308 119
rect 1313 116 1341 119
rect 1346 116 1349 119
rect 977 110 980 113
rect 985 110 1013 113
rect 1018 110 1021 113
rect 1108 106 1111 109
rect 1116 106 1144 109
rect 1149 106 1152 109
rect 1305 106 1308 109
rect 1313 106 1316 109
rect 977 100 980 103
rect 985 100 988 103
rect 993 100 1013 103
rect 1018 100 1021 103
rect 1321 106 1341 109
rect 1346 106 1349 109
rect 1735 124 1738 127
rect 1746 124 1749 127
rect 1517 121 1532 124
rect 1540 121 1543 124
rect 1576 121 1579 124
rect 1587 121 1601 124
rect 1605 121 1611 124
rect 1619 121 1622 124
rect 1434 104 1447 107
rect 1455 104 1479 107
rect 1487 104 1490 107
rect 1497 104 1500 107
rect 1508 104 1532 107
rect 1540 104 1552 107
rect 1108 96 1111 99
rect 1116 96 1144 99
rect 1149 96 1152 99
rect 1108 86 1111 89
rect 1116 86 1119 89
rect 1124 86 1144 89
rect 1149 86 1152 89
rect 1567 104 1579 107
rect 1587 104 1611 107
rect 1619 104 1622 107
rect 1755 124 1770 127
rect 1778 124 1781 127
rect 1814 124 1817 127
rect 1825 124 1839 127
rect 1843 124 1849 127
rect 1857 124 1860 127
rect 1968 124 1971 127
rect 1979 124 1982 127
rect 1672 107 1685 110
rect 1693 107 1717 110
rect 1725 107 1728 110
rect 1735 107 1738 110
rect 1746 107 1770 110
rect 1778 107 1790 110
rect 1434 87 1447 90
rect 1455 87 1479 90
rect 1487 87 1490 90
rect 1805 107 1817 110
rect 1825 107 1849 110
rect 1857 107 1860 110
rect 2206 127 2209 130
rect 2217 127 2220 130
rect 1988 124 2003 127
rect 2011 124 2014 127
rect 2047 124 2050 127
rect 2058 124 2072 127
rect 2076 124 2082 127
rect 2090 124 2093 127
rect 1905 107 1918 110
rect 1926 107 1950 110
rect 1958 107 1961 110
rect 1968 107 1971 110
rect 1979 107 2003 110
rect 2011 107 2023 110
rect 1672 90 1685 93
rect 1693 90 1717 93
rect 1725 90 1728 93
rect 764 78 767 81
rect 772 78 800 81
rect 805 78 808 81
rect 2038 107 2050 110
rect 2058 107 2082 110
rect 2090 107 2093 110
rect 2226 127 2241 130
rect 2249 127 2252 130
rect 2285 127 2288 130
rect 2296 127 2310 130
rect 2314 127 2320 130
rect 2328 127 2331 130
rect 2143 110 2156 113
rect 2164 110 2188 113
rect 2196 110 2199 113
rect 2206 110 2209 113
rect 2217 110 2241 113
rect 2249 110 2261 113
rect 1905 90 1918 93
rect 1926 90 1950 93
rect 1958 90 1961 93
rect 2454 126 2457 141
rect 2454 117 2457 121
rect 2504 117 2507 141
rect 2521 117 2524 141
rect 2276 110 2288 113
rect 2296 110 2320 113
rect 2328 110 2331 113
rect 2454 106 2457 109
rect 2504 99 2507 109
rect 2521 99 2524 109
rect 2143 93 2156 96
rect 2164 93 2188 96
rect 2196 93 2199 96
rect 2373 93 2376 96
rect 2384 93 2408 96
rect 2416 93 2426 96
rect 764 68 767 71
rect 772 68 800 71
rect 805 68 808 71
rect 2258 74 2261 77
rect 2275 74 2278 77
rect 2373 76 2376 79
rect 2384 76 2408 79
rect 2416 76 2426 79
rect 1787 71 1790 74
rect 1804 71 1807 74
rect 2020 71 2023 74
rect 2037 71 2040 74
rect 1300 65 1303 68
rect 1311 65 1317 68
rect 764 58 767 61
rect 772 58 775 61
rect 780 58 800 61
rect 805 58 808 61
rect 972 59 975 62
rect 983 59 989 62
rect 1549 68 1552 71
rect 1566 68 1569 71
rect 1322 65 1335 68
rect 1343 65 1346 68
rect 994 59 1007 62
rect 1015 59 1018 62
rect 1103 45 1106 48
rect 1114 45 1120 48
rect 1125 45 1138 48
rect 1146 45 1149 48
rect 1549 35 1552 60
rect 1566 35 1569 60
rect 1787 38 1790 63
rect 1804 38 1807 63
rect 2020 38 2023 63
rect 2037 38 2040 63
rect 2258 41 2261 66
rect 2275 41 2278 66
rect 2454 61 2457 64
rect 2504 61 2507 71
rect 2521 61 2524 71
rect 2454 49 2457 53
rect 2258 30 2261 33
rect 2275 30 2278 33
rect 1787 27 1790 30
rect 1804 27 1807 30
rect 2020 27 2023 30
rect 2037 27 2040 30
rect 1549 24 1552 27
rect 1566 24 1569 27
rect 759 17 762 20
rect 770 17 776 20
rect 781 17 794 20
rect 802 17 805 20
rect 1431 13 1434 16
rect 1442 13 1457 16
rect 1669 16 1672 19
rect 1680 16 1695 19
rect 1462 13 1466 16
rect 1474 13 1477 16
rect 1700 16 1704 19
rect 1712 16 1715 19
rect 1902 16 1905 19
rect 1913 16 1928 19
rect 2454 29 2457 44
rect 2504 29 2507 53
rect 2521 29 2524 53
rect 2140 19 2143 22
rect 2151 19 2166 22
rect 1933 16 1937 19
rect 1945 16 1948 19
rect 2171 19 2175 22
rect 2183 19 2186 22
rect 2454 18 2457 21
rect 2504 18 2507 21
rect 2521 18 2524 21
rect 1135 -10 1138 -7
rect 1146 -10 1152 -7
rect 819 -24 822 -21
rect 830 -24 836 -21
rect 907 -19 910 -16
rect 918 -19 924 -16
rect 841 -24 854 -21
rect 862 -24 865 -21
rect 1157 -10 1170 -7
rect 1178 -10 1181 -7
rect 929 -19 942 -16
rect 950 -19 953 -16
rect 1237 -12 1240 -9
rect 1248 -12 1254 -9
rect 1259 -12 1272 -9
rect 1280 -12 1283 -9
rect 2373 -16 2376 -13
rect 2384 -16 2399 -13
rect 2454 -10 2457 -7
rect 2504 -10 2507 -7
rect 2521 -10 2524 -7
rect 2404 -16 2408 -13
rect 2416 -16 2419 -13
rect 2259 -22 2262 -19
rect 2276 -22 2279 -19
rect 1788 -25 1791 -22
rect 1805 -25 1808 -22
rect 2021 -25 2024 -22
rect 2038 -25 2041 -22
rect 1550 -28 1553 -25
rect 1567 -28 1570 -25
rect 1136 -45 1139 -42
rect 1144 -45 1172 -42
rect 1177 -45 1180 -42
rect 908 -54 911 -51
rect 916 -54 944 -51
rect 949 -54 952 -51
rect 820 -59 823 -56
rect 828 -59 856 -56
rect 861 -59 864 -56
rect 1238 -47 1241 -44
rect 1246 -47 1274 -44
rect 1279 -47 1282 -44
rect 1136 -55 1139 -52
rect 1144 -55 1172 -52
rect 1177 -55 1180 -52
rect 908 -64 911 -61
rect 916 -64 944 -61
rect 949 -64 952 -61
rect 1238 -57 1241 -54
rect 1246 -57 1274 -54
rect 1279 -57 1282 -54
rect 1431 -55 1434 -52
rect 1442 -55 1466 -52
rect 1474 -55 1484 -52
rect 820 -69 823 -66
rect 828 -69 856 -66
rect 861 -69 864 -66
rect 1136 -65 1139 -62
rect 1144 -65 1147 -62
rect 908 -74 911 -71
rect 916 -74 919 -71
rect 820 -79 823 -76
rect 828 -79 831 -76
rect 1152 -65 1172 -62
rect 1177 -65 1180 -62
rect 1238 -67 1241 -64
rect 1246 -67 1249 -64
rect 1254 -67 1274 -64
rect 1279 -67 1282 -64
rect 924 -74 944 -71
rect 949 -74 952 -71
rect 1550 -60 1553 -36
rect 1567 -60 1570 -36
rect 1669 -52 1672 -49
rect 1680 -52 1704 -49
rect 1712 -52 1722 -49
rect 1788 -57 1791 -33
rect 1805 -57 1808 -33
rect 1902 -52 1905 -49
rect 1913 -52 1937 -49
rect 1945 -52 1955 -49
rect 1431 -72 1434 -69
rect 1442 -72 1466 -69
rect 1474 -72 1484 -69
rect 836 -79 856 -76
rect 861 -79 864 -76
rect 1550 -71 1553 -68
rect 1567 -71 1570 -68
rect 1669 -69 1672 -66
rect 1680 -69 1704 -66
rect 1712 -69 1722 -66
rect 1788 -68 1791 -65
rect 1805 -68 1808 -65
rect 2021 -57 2024 -33
rect 2038 -57 2041 -33
rect 2140 -49 2143 -46
rect 2151 -49 2175 -46
rect 2183 -49 2193 -46
rect 2259 -54 2262 -30
rect 2276 -54 2279 -30
rect 2454 -33 2457 -18
rect 2454 -42 2457 -38
rect 2504 -42 2507 -18
rect 2521 -42 2524 -18
rect 2454 -53 2457 -50
rect 1902 -69 1905 -66
rect 1913 -69 1937 -66
rect 1945 -69 1955 -66
rect 2021 -68 2024 -65
rect 2038 -68 2041 -65
rect 2140 -66 2143 -63
rect 2151 -66 2175 -63
rect 2183 -66 2193 -63
rect 2259 -65 2262 -62
rect 2276 -65 2279 -62
rect 2504 -60 2507 -50
rect 2521 -60 2524 -50
rect 2373 -66 2376 -63
rect 2384 -66 2408 -63
rect 2416 -66 2426 -63
rect 2373 -83 2376 -80
rect 2384 -83 2408 -80
rect 2416 -83 2426 -80
rect 1131 -106 1134 -103
rect 1142 -106 1148 -103
rect 815 -120 818 -117
rect 826 -120 832 -117
rect 903 -115 906 -112
rect 914 -115 920 -112
rect 837 -120 850 -117
rect 858 -120 861 -117
rect 1153 -106 1166 -103
rect 1174 -106 1177 -103
rect 925 -115 938 -112
rect 946 -115 949 -112
rect 1233 -108 1236 -105
rect 1244 -108 1250 -105
rect 1497 -103 1500 -100
rect 1508 -103 1511 -100
rect 1255 -108 1268 -105
rect 1276 -108 1279 -105
rect 1735 -100 1738 -97
rect 1746 -100 1749 -97
rect 1517 -103 1532 -100
rect 1540 -103 1543 -100
rect 1576 -103 1579 -100
rect 1587 -103 1601 -100
rect 1605 -103 1611 -100
rect 1619 -103 1622 -100
rect 1497 -120 1500 -117
rect 1508 -120 1532 -117
rect 1540 -120 1552 -117
rect 1432 -128 1435 -125
rect 1443 -128 1458 -125
rect 1463 -128 1467 -125
rect 1475 -128 1478 -125
rect 1755 -100 1770 -97
rect 1778 -100 1781 -97
rect 1814 -100 1817 -97
rect 1825 -100 1839 -97
rect 1843 -100 1849 -97
rect 1857 -100 1860 -97
rect 1968 -100 1971 -97
rect 1979 -100 1982 -97
rect 1567 -120 1579 -117
rect 1587 -120 1611 -117
rect 1619 -120 1622 -117
rect 1735 -117 1738 -114
rect 1746 -117 1770 -114
rect 1778 -117 1790 -114
rect 1670 -125 1673 -122
rect 1681 -125 1696 -122
rect 1701 -125 1705 -122
rect 1713 -125 1716 -122
rect 2206 -97 2209 -94
rect 2217 -97 2220 -94
rect 1988 -100 2003 -97
rect 2011 -100 2014 -97
rect 2047 -100 2050 -97
rect 2058 -100 2072 -97
rect 2076 -100 2082 -97
rect 2090 -100 2093 -97
rect 1805 -117 1817 -114
rect 1825 -117 1849 -114
rect 1857 -117 1860 -114
rect 1968 -117 1971 -114
rect 1979 -117 2003 -114
rect 2011 -117 2023 -114
rect 1903 -125 1906 -122
rect 1914 -125 1929 -122
rect 1934 -125 1938 -122
rect 1946 -125 1949 -122
rect 2226 -97 2241 -94
rect 2249 -97 2252 -94
rect 2285 -97 2288 -94
rect 2296 -97 2310 -94
rect 2314 -97 2320 -94
rect 2328 -97 2331 -94
rect 2038 -117 2050 -114
rect 2058 -117 2082 -114
rect 2090 -117 2093 -114
rect 2206 -114 2209 -111
rect 2217 -114 2241 -111
rect 2249 -114 2261 -111
rect 2141 -122 2144 -119
rect 2152 -122 2167 -119
rect 2172 -122 2176 -119
rect 2184 -122 2187 -119
rect 2454 -98 2457 -95
rect 2504 -98 2507 -88
rect 2521 -98 2524 -88
rect 2454 -110 2457 -106
rect 2276 -114 2288 -111
rect 2296 -114 2320 -111
rect 2328 -114 2331 -111
rect 2454 -130 2457 -115
rect 2504 -130 2507 -106
rect 2521 -130 2524 -106
rect 2454 -141 2457 -138
rect 2504 -141 2507 -138
rect 2521 -141 2524 -138
rect 2258 -150 2261 -147
rect 2275 -150 2278 -147
rect 1787 -153 1790 -150
rect 1804 -153 1807 -150
rect 2020 -153 2023 -150
rect 2037 -153 2040 -150
rect 1549 -156 1552 -153
rect 1566 -156 1569 -153
rect 1353 -183 1356 -180
rect 1364 -183 1368 -180
rect 1373 -183 1388 -180
rect 1396 -183 1399 -180
rect 972 -200 975 -197
rect 983 -200 987 -197
rect 992 -200 1007 -197
rect 1015 -200 1018 -197
rect 1122 -200 1125 -197
rect 1133 -200 1137 -197
rect 1549 -189 1552 -164
rect 1566 -189 1569 -164
rect 1142 -200 1157 -197
rect 1165 -200 1168 -197
rect 1269 -200 1272 -197
rect 1280 -200 1284 -197
rect 1432 -196 1435 -193
rect 1443 -196 1467 -193
rect 1475 -196 1485 -193
rect 1289 -200 1304 -197
rect 1312 -200 1315 -197
rect 1787 -186 1790 -161
rect 1804 -186 1807 -161
rect 1670 -193 1673 -190
rect 1681 -193 1705 -190
rect 1713 -193 1723 -190
rect 1549 -200 1552 -197
rect 1566 -200 1569 -197
rect 2020 -186 2023 -161
rect 2037 -186 2040 -161
rect 1903 -193 1906 -190
rect 1914 -193 1938 -190
rect 1946 -193 1956 -190
rect 1787 -197 1790 -194
rect 1804 -197 1807 -194
rect 1432 -213 1435 -210
rect 1443 -213 1467 -210
rect 1475 -213 1485 -210
rect 1670 -210 1673 -207
rect 1681 -210 1705 -207
rect 1713 -210 1723 -207
rect 2258 -183 2261 -158
rect 2275 -183 2278 -158
rect 2372 -170 2375 -167
rect 2383 -170 2398 -167
rect 2453 -164 2456 -161
rect 2503 -164 2506 -161
rect 2520 -164 2523 -161
rect 2403 -170 2407 -167
rect 2415 -170 2418 -167
rect 2141 -190 2144 -187
rect 2152 -190 2176 -187
rect 2184 -190 2194 -187
rect 2020 -197 2023 -194
rect 2037 -197 2040 -194
rect 2453 -187 2456 -172
rect 2258 -194 2261 -191
rect 2275 -194 2278 -191
rect 2453 -196 2456 -192
rect 2503 -196 2506 -172
rect 2520 -196 2523 -172
rect 1903 -210 1906 -207
rect 1914 -210 1938 -207
rect 1946 -210 1956 -207
rect 2141 -207 2144 -204
rect 2152 -207 2176 -204
rect 2184 -207 2194 -204
rect 2453 -207 2456 -204
rect 2503 -214 2506 -204
rect 2520 -214 2523 -204
rect 2372 -220 2375 -217
rect 2383 -220 2407 -217
rect 2415 -220 2425 -217
rect 1346 -233 1356 -230
rect 1364 -233 1388 -230
rect 1396 -233 1399 -230
rect 965 -250 975 -247
rect 983 -250 1007 -247
rect 1015 -250 1018 -247
rect 569 -272 572 -269
rect 577 -272 585 -269
rect 1115 -250 1125 -247
rect 1133 -250 1157 -247
rect 1165 -250 1168 -247
rect 965 -267 975 -264
rect 983 -267 1007 -264
rect 1015 -267 1018 -264
rect 590 -272 605 -269
rect 610 -272 613 -269
rect 1262 -250 1272 -247
rect 1280 -250 1304 -247
rect 1312 -250 1315 -247
rect 1115 -267 1125 -264
rect 1133 -267 1157 -264
rect 1165 -267 1168 -264
rect 2372 -237 2375 -234
rect 2383 -237 2407 -234
rect 2415 -237 2425 -234
rect 1346 -250 1356 -247
rect 1364 -250 1388 -247
rect 1396 -250 1399 -247
rect 2182 -254 2185 -251
rect 2199 -254 2202 -251
rect 2453 -252 2456 -249
rect 2503 -252 2506 -242
rect 2520 -252 2523 -242
rect 1711 -257 1714 -254
rect 1728 -257 1731 -254
rect 1944 -257 1947 -254
rect 1961 -257 1964 -254
rect 1473 -260 1476 -257
rect 1490 -260 1493 -257
rect 1262 -267 1272 -264
rect 1280 -267 1304 -264
rect 1312 -267 1315 -264
rect 757 -292 760 -289
rect 768 -292 774 -289
rect 779 -292 792 -289
rect 800 -292 803 -289
rect 913 -292 916 -289
rect 924 -292 930 -289
rect 935 -292 948 -289
rect 956 -292 959 -289
rect 1063 -292 1066 -289
rect 1074 -292 1080 -289
rect 1085 -292 1098 -289
rect 1106 -292 1109 -289
rect 1210 -292 1213 -289
rect 1221 -292 1227 -289
rect 1232 -292 1245 -289
rect 1253 -292 1256 -289
rect 1473 -292 1476 -268
rect 1490 -292 1493 -268
rect 1711 -289 1714 -265
rect 1728 -289 1731 -265
rect 1944 -289 1947 -265
rect 1961 -289 1964 -265
rect 2182 -286 2185 -262
rect 2199 -286 2202 -262
rect 2453 -264 2456 -260
rect 2453 -284 2456 -269
rect 2503 -284 2506 -260
rect 2520 -284 2523 -260
rect 2182 -297 2185 -294
rect 2199 -297 2202 -294
rect 2453 -295 2456 -292
rect 2503 -295 2506 -292
rect 2520 -295 2523 -292
rect 1711 -300 1714 -297
rect 1728 -300 1731 -297
rect 1944 -300 1947 -297
rect 1961 -300 1964 -297
rect 1473 -303 1476 -300
rect 1490 -303 1493 -300
rect 569 -306 572 -303
rect 577 -306 605 -303
rect 610 -306 613 -303
rect 569 -316 572 -313
rect 577 -316 605 -313
rect 610 -316 613 -313
rect 803 -318 806 -315
rect 820 -318 823 -315
rect 959 -318 962 -315
rect 976 -318 979 -315
rect 1109 -318 1112 -315
rect 1126 -318 1129 -315
rect 1256 -318 1259 -315
rect 1273 -318 1276 -315
rect 569 -326 572 -323
rect 577 -326 605 -323
rect 610 -326 613 -323
rect 654 -348 667 -345
rect 675 -348 699 -345
rect 707 -348 710 -345
rect 803 -350 806 -326
rect 820 -350 823 -326
rect 959 -350 962 -326
rect 976 -350 979 -326
rect 1109 -350 1112 -326
rect 1126 -350 1129 -326
rect 1256 -350 1259 -326
rect 1273 -350 1276 -326
rect 1420 -335 1423 -332
rect 1431 -335 1434 -332
rect 1658 -332 1661 -329
rect 1669 -332 1672 -329
rect 1440 -335 1455 -332
rect 1463 -335 1466 -332
rect 1499 -335 1502 -332
rect 1510 -335 1524 -332
rect 1528 -335 1534 -332
rect 1542 -335 1545 -332
rect 1420 -352 1423 -349
rect 1431 -352 1455 -349
rect 1463 -352 1475 -349
rect 803 -361 806 -358
rect 820 -361 823 -358
rect 959 -361 962 -358
rect 976 -361 979 -358
rect 1109 -361 1112 -358
rect 1126 -361 1129 -358
rect 1256 -361 1259 -358
rect 1273 -361 1276 -358
rect 1678 -332 1693 -329
rect 1701 -332 1704 -329
rect 1737 -332 1740 -329
rect 1748 -332 1762 -329
rect 1766 -332 1772 -329
rect 1780 -332 1783 -329
rect 1891 -332 1894 -329
rect 1902 -332 1905 -329
rect 1658 -349 1661 -346
rect 1669 -349 1693 -346
rect 1701 -349 1713 -346
rect 1490 -352 1502 -349
rect 1510 -352 1534 -349
rect 1542 -352 1545 -349
rect 2129 -329 2132 -326
rect 2140 -329 2143 -326
rect 1911 -332 1926 -329
rect 1934 -332 1937 -329
rect 1970 -332 1973 -329
rect 1981 -332 1995 -329
rect 1999 -332 2005 -329
rect 2013 -332 2016 -329
rect 1728 -349 1740 -346
rect 1748 -349 1772 -346
rect 1780 -349 1783 -346
rect 1891 -349 1894 -346
rect 1902 -349 1926 -346
rect 1934 -349 1946 -346
rect 2149 -329 2164 -326
rect 2172 -329 2175 -326
rect 2208 -329 2211 -326
rect 2219 -329 2233 -326
rect 2237 -329 2243 -326
rect 2251 -329 2254 -326
rect 2372 -329 2375 -326
rect 2383 -329 2398 -326
rect 2129 -346 2132 -343
rect 2140 -346 2164 -343
rect 2172 -346 2184 -343
rect 1961 -349 1973 -346
rect 1981 -349 2005 -346
rect 2013 -349 2016 -346
rect 2453 -323 2456 -320
rect 2503 -323 2506 -320
rect 2520 -323 2523 -320
rect 2403 -329 2407 -326
rect 2415 -329 2418 -326
rect 2199 -346 2211 -343
rect 2219 -346 2243 -343
rect 2251 -346 2254 -343
rect 2453 -346 2456 -331
rect 2453 -355 2456 -351
rect 2503 -355 2506 -331
rect 2520 -355 2523 -331
rect 654 -365 667 -362
rect 675 -365 699 -362
rect 707 -365 710 -362
rect 2453 -366 2456 -363
rect 2503 -373 2506 -363
rect 2520 -373 2523 -363
rect 2372 -379 2375 -376
rect 2383 -379 2407 -376
rect 2415 -379 2425 -376
rect 569 -385 572 -382
rect 577 -385 585 -382
rect 2181 -382 2184 -379
rect 2198 -382 2201 -379
rect 590 -385 605 -382
rect 610 -385 613 -382
rect 750 -393 753 -390
rect 761 -393 764 -390
rect 664 -405 667 -402
rect 675 -405 690 -402
rect 695 -405 699 -402
rect 707 -405 710 -402
rect 770 -393 785 -390
rect 793 -393 796 -390
rect 829 -393 832 -390
rect 840 -393 854 -390
rect 858 -393 864 -390
rect 872 -393 875 -390
rect 906 -393 909 -390
rect 917 -393 920 -390
rect 750 -410 753 -407
rect 761 -410 785 -407
rect 793 -410 805 -407
rect 569 -419 572 -416
rect 577 -419 605 -416
rect 610 -419 613 -416
rect 926 -393 941 -390
rect 949 -393 952 -390
rect 985 -393 988 -390
rect 996 -393 1010 -390
rect 1014 -393 1020 -390
rect 1028 -393 1031 -390
rect 1056 -393 1059 -390
rect 1067 -393 1070 -390
rect 820 -410 832 -407
rect 840 -410 864 -407
rect 872 -410 875 -407
rect 906 -410 909 -407
rect 917 -410 941 -407
rect 949 -410 961 -407
rect 1076 -393 1091 -390
rect 1099 -393 1102 -390
rect 1135 -393 1138 -390
rect 1146 -393 1160 -390
rect 1164 -393 1170 -390
rect 1178 -393 1181 -390
rect 1203 -393 1206 -390
rect 1214 -393 1217 -390
rect 976 -410 988 -407
rect 996 -410 1020 -407
rect 1028 -410 1031 -407
rect 1056 -410 1059 -407
rect 1067 -410 1091 -407
rect 1099 -410 1111 -407
rect 1710 -385 1713 -382
rect 1727 -385 1730 -382
rect 1943 -385 1946 -382
rect 1960 -385 1963 -382
rect 1472 -388 1475 -385
rect 1489 -388 1492 -385
rect 1223 -393 1238 -390
rect 1246 -393 1249 -390
rect 1282 -393 1285 -390
rect 1293 -393 1307 -390
rect 1311 -393 1317 -390
rect 1325 -393 1328 -390
rect 1126 -410 1138 -407
rect 1146 -410 1170 -407
rect 1178 -410 1181 -407
rect 1203 -410 1206 -407
rect 1214 -410 1238 -407
rect 1246 -410 1258 -407
rect 1273 -410 1285 -407
rect 1293 -410 1317 -407
rect 1325 -410 1328 -407
rect 1472 -421 1475 -396
rect 1489 -421 1492 -396
rect 1710 -418 1713 -393
rect 1727 -418 1730 -393
rect 1943 -418 1946 -393
rect 1960 -418 1963 -393
rect 2181 -415 2184 -390
rect 2198 -415 2201 -390
rect 2372 -396 2375 -393
rect 2383 -396 2407 -393
rect 2415 -396 2425 -393
rect 2453 -411 2456 -408
rect 2503 -411 2506 -401
rect 2520 -411 2523 -401
rect 569 -429 572 -426
rect 577 -429 605 -426
rect 610 -429 613 -426
rect 2453 -423 2456 -419
rect 2181 -426 2184 -423
rect 2198 -426 2201 -423
rect 1710 -429 1713 -426
rect 1727 -429 1730 -426
rect 1943 -429 1946 -426
rect 1960 -429 1963 -426
rect 1472 -432 1475 -429
rect 1489 -432 1492 -429
rect 569 -439 572 -436
rect 577 -439 605 -436
rect 610 -439 613 -436
rect 2453 -443 2456 -428
rect 2503 -443 2506 -419
rect 2520 -443 2523 -419
rect 802 -446 805 -443
rect 819 -446 822 -443
rect 958 -446 961 -443
rect 975 -446 978 -443
rect 1108 -446 1111 -443
rect 1125 -446 1128 -443
rect 1255 -446 1258 -443
rect 1272 -446 1275 -443
rect 2453 -454 2456 -451
rect 2503 -454 2506 -451
rect 2520 -454 2523 -451
rect 462 -483 465 -480
rect 470 -483 485 -480
rect 802 -479 805 -454
rect 819 -479 822 -454
rect 958 -479 961 -454
rect 975 -479 978 -454
rect 1108 -479 1111 -454
rect 1125 -479 1128 -454
rect 1255 -479 1258 -454
rect 1272 -479 1275 -454
rect 490 -483 498 -480
rect 503 -483 506 -480
rect 569 -493 572 -490
rect 577 -493 585 -490
rect 802 -490 805 -487
rect 819 -490 822 -487
rect 958 -490 961 -487
rect 975 -490 978 -487
rect 1108 -490 1111 -487
rect 1125 -490 1128 -487
rect 1255 -490 1258 -487
rect 1272 -490 1275 -487
rect 590 -493 605 -490
rect 610 -493 613 -490
rect 753 -523 756 -520
rect 764 -523 779 -520
rect 569 -527 572 -524
rect 577 -527 605 -524
rect 610 -527 613 -524
rect 784 -523 788 -520
rect 796 -523 799 -520
rect 835 -523 838 -520
rect 846 -523 850 -520
rect 855 -523 870 -520
rect 878 -523 881 -520
rect 909 -523 912 -520
rect 920 -523 935 -520
rect 940 -523 944 -520
rect 952 -523 955 -520
rect 991 -523 994 -520
rect 1002 -523 1006 -520
rect 1011 -523 1026 -520
rect 1034 -523 1037 -520
rect 1059 -523 1062 -520
rect 1070 -523 1085 -520
rect 1090 -523 1094 -520
rect 1102 -523 1105 -520
rect 1141 -523 1144 -520
rect 1152 -523 1156 -520
rect 1161 -523 1176 -520
rect 1184 -523 1187 -520
rect 1215 -523 1218 -520
rect 1226 -523 1241 -520
rect 1246 -523 1250 -520
rect 1258 -523 1261 -520
rect 1297 -523 1300 -520
rect 1308 -523 1312 -520
rect 1317 -523 1332 -520
rect 1340 -523 1343 -520
rect 1461 -523 1464 -520
rect 1472 -523 1487 -520
rect 1492 -523 1496 -520
rect 1504 -523 1507 -520
rect 1550 -523 1553 -520
rect 1561 -523 1565 -520
rect 1570 -523 1585 -520
rect 1593 -523 1596 -520
rect 1700 -522 1703 -519
rect 1711 -522 1726 -519
rect 1731 -522 1735 -519
rect 1743 -522 1746 -519
rect 1788 -522 1791 -519
rect 1799 -522 1803 -519
rect 1808 -522 1823 -519
rect 1831 -522 1834 -519
rect 1933 -522 1936 -519
rect 1944 -522 1959 -519
rect 1964 -522 1968 -519
rect 1976 -522 1979 -519
rect 2021 -522 2024 -519
rect 2032 -522 2036 -519
rect 2041 -522 2056 -519
rect 2064 -522 2067 -519
rect 2154 -522 2157 -519
rect 2165 -522 2180 -519
rect 2185 -522 2189 -519
rect 2197 -522 2200 -519
rect 2242 -522 2245 -519
rect 2253 -522 2257 -519
rect 2262 -522 2277 -519
rect 2285 -522 2288 -519
rect 2324 -525 2327 -522
rect 2335 -525 2339 -522
rect 2344 -525 2359 -522
rect 2367 -525 2370 -522
rect 569 -537 572 -534
rect 577 -537 605 -534
rect 610 -537 613 -534
rect 569 -547 572 -544
rect 577 -547 605 -544
rect 610 -547 613 -544
rect 1461 -578 1464 -575
rect 1472 -578 1496 -575
rect 1504 -578 1514 -575
rect 427 -589 430 -586
rect 435 -589 443 -586
rect 448 -589 463 -586
rect 468 -589 471 -586
rect 753 -588 756 -585
rect 764 -588 788 -585
rect 796 -588 806 -585
rect 569 -604 572 -601
rect 577 -604 585 -601
rect 590 -604 605 -601
rect 610 -604 613 -601
rect 828 -588 838 -585
rect 846 -588 870 -585
rect 878 -588 881 -585
rect 909 -588 912 -585
rect 920 -588 944 -585
rect 952 -588 962 -585
rect 753 -605 756 -602
rect 764 -605 788 -602
rect 796 -605 806 -602
rect 984 -588 994 -585
rect 1002 -588 1026 -585
rect 1034 -588 1037 -585
rect 1059 -588 1062 -585
rect 1070 -588 1094 -585
rect 1102 -588 1112 -585
rect 828 -605 838 -602
rect 846 -605 870 -602
rect 878 -605 881 -602
rect 909 -605 912 -602
rect 920 -605 944 -602
rect 952 -605 962 -602
rect 1134 -588 1144 -585
rect 1152 -588 1176 -585
rect 1184 -588 1187 -585
rect 1215 -588 1218 -585
rect 1226 -588 1250 -585
rect 1258 -588 1268 -585
rect 984 -605 994 -602
rect 1002 -605 1026 -602
rect 1034 -605 1037 -602
rect 1059 -605 1062 -602
rect 1070 -605 1094 -602
rect 1102 -605 1112 -602
rect 1290 -588 1300 -585
rect 1308 -588 1332 -585
rect 1340 -588 1343 -585
rect 1134 -605 1144 -602
rect 1152 -605 1176 -602
rect 1184 -605 1187 -602
rect 1215 -605 1218 -602
rect 1226 -605 1250 -602
rect 1258 -605 1268 -602
rect 1543 -578 1553 -575
rect 1561 -578 1585 -575
rect 1593 -578 1596 -575
rect 1700 -577 1703 -574
rect 1711 -577 1735 -574
rect 1743 -577 1753 -574
rect 1461 -595 1464 -592
rect 1472 -595 1496 -592
rect 1504 -595 1514 -592
rect 1290 -605 1300 -602
rect 1308 -605 1332 -602
rect 1340 -605 1343 -602
rect 1781 -577 1791 -574
rect 1799 -577 1823 -574
rect 1831 -577 1834 -574
rect 1933 -577 1936 -574
rect 1944 -577 1968 -574
rect 1976 -577 1986 -574
rect 1543 -595 1553 -592
rect 1561 -595 1585 -592
rect 1593 -595 1596 -592
rect 1700 -594 1703 -591
rect 1711 -594 1735 -591
rect 1743 -594 1753 -591
rect 2014 -577 2024 -574
rect 2032 -577 2056 -574
rect 2064 -577 2067 -574
rect 2154 -577 2157 -574
rect 2165 -577 2189 -574
rect 2197 -577 2207 -574
rect 1781 -594 1791 -591
rect 1799 -594 1823 -591
rect 1831 -594 1834 -591
rect 1933 -594 1936 -591
rect 1944 -594 1968 -591
rect 1976 -594 1986 -591
rect 2235 -577 2245 -574
rect 2253 -577 2277 -574
rect 2285 -577 2288 -574
rect 2014 -594 2024 -591
rect 2032 -594 2056 -591
rect 2064 -594 2067 -591
rect 2154 -594 2157 -591
rect 2165 -594 2189 -591
rect 2197 -594 2207 -591
rect 2317 -580 2327 -577
rect 2335 -580 2359 -577
rect 2367 -580 2370 -577
rect 2235 -594 2245 -591
rect 2253 -594 2277 -591
rect 2285 -594 2288 -591
rect 2317 -597 2327 -594
rect 2335 -597 2359 -594
rect 2367 -597 2370 -594
rect 569 -638 572 -635
rect 577 -638 605 -635
rect 610 -638 613 -635
rect 569 -648 572 -645
rect 577 -648 605 -645
rect 610 -648 613 -645
rect 569 -658 572 -655
rect 577 -658 605 -655
rect 610 -658 613 -655
<< polycontact >>
rect 1614 327 1619 332
rect 1751 322 1756 327
rect 1895 324 1900 329
rect 2038 325 2043 330
rect 1694 291 1699 296
rect 1704 291 1709 296
rect 1714 291 1719 296
rect 1838 293 1843 298
rect 1848 293 1853 298
rect 1858 293 1863 298
rect 1981 294 1986 299
rect 1991 294 1996 299
rect 2001 294 2006 299
rect 1557 287 1562 291
rect 1574 287 1579 291
rect 1032 240 1037 245
rect 1101 240 1106 245
rect 968 209 973 214
rect 978 209 983 214
rect 988 209 993 214
rect 998 209 1003 214
rect 1135 209 1140 214
rect 1145 209 1150 214
rect 1155 209 1160 214
rect 1165 209 1170 214
rect 993 154 998 159
rect 1321 160 1326 165
rect 1124 140 1129 145
rect 1470 143 1475 148
rect 1549 149 1554 153
rect 1566 149 1571 153
rect 1708 146 1713 151
rect 1787 152 1792 156
rect 1804 152 1809 156
rect 1941 146 1946 151
rect 2020 152 2025 156
rect 2037 152 2042 156
rect 2179 149 2184 154
rect 2258 155 2263 159
rect 2275 155 2280 159
rect 2399 142 2404 147
rect 972 119 977 124
rect 1300 125 1305 130
rect 780 112 785 117
rect 972 109 977 114
rect 1300 115 1305 120
rect 1103 105 1108 110
rect 988 99 993 104
rect 1103 95 1108 100
rect 1316 105 1321 110
rect 1430 103 1434 108
rect 1511 120 1517 125
rect 1601 120 1605 124
rect 759 77 764 82
rect 1119 85 1124 90
rect 1430 86 1434 91
rect 1552 103 1557 108
rect 1562 103 1567 108
rect 1668 106 1672 111
rect 1749 123 1755 128
rect 1839 123 1843 127
rect 1668 89 1672 94
rect 1790 106 1795 111
rect 1800 106 1805 111
rect 1901 106 1905 111
rect 1982 123 1988 128
rect 2072 123 2076 127
rect 1901 89 1905 94
rect 2023 106 2028 111
rect 2033 106 2038 111
rect 2139 109 2143 114
rect 2220 126 2226 131
rect 2310 126 2314 130
rect 2139 92 2143 97
rect 2261 109 2266 114
rect 2271 109 2276 114
rect 2453 121 2458 126
rect 2426 92 2430 97
rect 2503 95 2508 99
rect 2520 95 2525 99
rect 759 67 764 72
rect 775 57 780 62
rect 989 58 994 63
rect 1317 64 1322 69
rect 2426 75 2430 80
rect 2503 71 2508 75
rect 2520 71 2525 75
rect 1120 44 1125 49
rect 2453 44 2458 49
rect 776 16 781 21
rect 1548 20 1553 24
rect 1565 20 1570 24
rect 1457 12 1462 17
rect 1786 23 1791 27
rect 1803 23 1808 27
rect 1695 15 1700 20
rect 2019 23 2024 27
rect 2036 23 2041 27
rect 1928 15 1933 20
rect 2257 26 2262 30
rect 2274 26 2279 30
rect 2166 18 2171 23
rect 836 -25 841 -20
rect 924 -20 929 -15
rect 1152 -11 1157 -6
rect 1254 -13 1259 -8
rect 2399 -17 2404 -12
rect 1131 -46 1136 -41
rect 815 -60 820 -55
rect 903 -55 908 -50
rect 815 -70 820 -65
rect 903 -65 908 -60
rect 1131 -56 1136 -51
rect 1233 -48 1238 -43
rect 1233 -58 1238 -53
rect 831 -80 836 -75
rect 919 -75 924 -70
rect 1147 -66 1152 -61
rect 1249 -68 1254 -63
rect 1484 -56 1488 -51
rect 1722 -53 1726 -48
rect 1484 -73 1488 -68
rect 1549 -75 1554 -71
rect 1566 -75 1571 -71
rect 1722 -70 1726 -65
rect 1955 -53 1959 -48
rect 2193 -50 2197 -45
rect 2453 -38 2458 -33
rect 1787 -72 1792 -68
rect 1804 -72 1809 -68
rect 1955 -70 1959 -65
rect 2020 -72 2025 -68
rect 2037 -72 2042 -68
rect 2193 -67 2197 -62
rect 2258 -69 2263 -65
rect 2275 -69 2280 -65
rect 2426 -67 2430 -62
rect 2503 -64 2508 -60
rect 2520 -64 2525 -60
rect 832 -121 837 -116
rect 920 -116 925 -111
rect 1148 -107 1153 -102
rect 1250 -109 1255 -104
rect 1511 -104 1517 -99
rect 1601 -104 1605 -100
rect 1458 -129 1463 -124
rect 1552 -121 1557 -116
rect 1562 -121 1567 -116
rect 1749 -101 1755 -96
rect 1839 -101 1843 -97
rect 1696 -126 1701 -121
rect 1790 -118 1795 -113
rect 1800 -118 1805 -113
rect 1982 -101 1988 -96
rect 2072 -101 2076 -97
rect 1929 -126 1934 -121
rect 2023 -118 2028 -113
rect 2033 -118 2038 -113
rect 2220 -98 2226 -93
rect 2426 -84 2430 -79
rect 2503 -88 2508 -84
rect 2520 -88 2525 -84
rect 2310 -98 2314 -94
rect 2167 -123 2172 -118
rect 2261 -115 2266 -110
rect 2271 -115 2276 -110
rect 2453 -115 2458 -110
rect 1368 -184 1373 -179
rect 987 -201 992 -196
rect 1137 -201 1142 -196
rect 1284 -201 1289 -196
rect 1485 -197 1489 -192
rect 1548 -204 1553 -200
rect 1565 -204 1570 -200
rect 1723 -194 1727 -189
rect 1786 -201 1791 -197
rect 1803 -201 1808 -197
rect 1485 -214 1489 -209
rect 1723 -211 1727 -206
rect 1956 -194 1960 -189
rect 2398 -171 2403 -166
rect 2019 -201 2024 -197
rect 2036 -201 2041 -197
rect 2194 -191 2198 -186
rect 2452 -192 2457 -187
rect 2257 -198 2262 -194
rect 2274 -198 2279 -194
rect 1956 -211 1960 -206
rect 2194 -208 2198 -203
rect 1342 -234 1346 -229
rect 961 -251 965 -246
rect 585 -273 590 -268
rect 961 -268 965 -263
rect 1111 -251 1115 -246
rect 1111 -268 1115 -263
rect 1258 -251 1262 -246
rect 1258 -268 1262 -263
rect 1342 -251 1346 -246
rect 2425 -221 2429 -216
rect 2502 -218 2507 -214
rect 2519 -218 2524 -214
rect 2425 -238 2429 -233
rect 2502 -242 2507 -238
rect 2519 -242 2524 -238
rect 774 -293 779 -288
rect 564 -307 569 -302
rect 930 -293 935 -288
rect 1080 -293 1085 -288
rect 1227 -293 1232 -288
rect 2452 -269 2457 -264
rect 564 -317 569 -312
rect 1472 -307 1477 -303
rect 1489 -307 1494 -303
rect 1710 -304 1715 -300
rect 1727 -304 1732 -300
rect 1943 -304 1948 -300
rect 1960 -304 1965 -300
rect 2181 -301 2186 -297
rect 2198 -301 2203 -297
rect 564 -327 569 -322
rect 650 -349 654 -344
rect 650 -366 654 -361
rect 1434 -336 1440 -331
rect 1524 -336 1528 -332
rect 1475 -353 1480 -348
rect 1485 -353 1490 -348
rect 1672 -333 1678 -328
rect 1762 -333 1766 -329
rect 1713 -350 1718 -345
rect 1723 -350 1728 -345
rect 1905 -333 1911 -328
rect 1995 -333 1999 -329
rect 1946 -350 1951 -345
rect 1956 -350 1961 -345
rect 2143 -330 2149 -325
rect 2233 -330 2237 -326
rect 2184 -347 2189 -342
rect 2194 -347 2199 -342
rect 2398 -330 2403 -325
rect 2452 -351 2457 -346
rect 802 -365 807 -361
rect 819 -365 824 -361
rect 958 -365 963 -361
rect 975 -365 980 -361
rect 1108 -365 1113 -361
rect 1125 -365 1130 -361
rect 1255 -365 1260 -361
rect 1272 -365 1277 -361
rect 585 -386 590 -381
rect 690 -406 695 -401
rect 564 -420 569 -415
rect 764 -394 770 -389
rect 854 -394 858 -390
rect 805 -411 810 -406
rect 815 -411 820 -406
rect 920 -394 926 -389
rect 1010 -394 1014 -390
rect 961 -411 966 -406
rect 971 -411 976 -406
rect 1070 -394 1076 -389
rect 1160 -394 1164 -390
rect 1111 -411 1116 -406
rect 1121 -411 1126 -406
rect 1217 -394 1223 -389
rect 1307 -394 1311 -390
rect 1258 -411 1263 -406
rect 1268 -411 1273 -406
rect 564 -430 569 -425
rect 2425 -380 2429 -375
rect 2502 -377 2507 -373
rect 2519 -377 2524 -373
rect 2425 -397 2429 -392
rect 2502 -401 2507 -397
rect 2519 -401 2524 -397
rect 564 -440 569 -435
rect 1471 -436 1476 -432
rect 1488 -436 1493 -432
rect 1709 -433 1714 -429
rect 1726 -433 1731 -429
rect 1942 -433 1947 -429
rect 1959 -433 1964 -429
rect 2180 -430 2185 -426
rect 2197 -430 2202 -426
rect 2452 -428 2457 -423
rect 485 -484 490 -479
rect 585 -494 590 -489
rect 801 -494 806 -490
rect 818 -494 823 -490
rect 957 -494 962 -490
rect 974 -494 979 -490
rect 1107 -494 1112 -490
rect 1124 -494 1129 -490
rect 1254 -494 1259 -490
rect 1271 -494 1276 -490
rect 564 -528 569 -523
rect 779 -524 784 -519
rect 564 -538 569 -533
rect 850 -524 855 -519
rect 935 -524 940 -519
rect 1006 -524 1011 -519
rect 1085 -524 1090 -519
rect 1156 -524 1161 -519
rect 1241 -524 1246 -519
rect 1312 -524 1317 -519
rect 1487 -524 1492 -519
rect 1565 -524 1570 -519
rect 1726 -523 1731 -518
rect 1803 -523 1808 -518
rect 1959 -523 1964 -518
rect 2036 -523 2041 -518
rect 2180 -523 2185 -518
rect 2257 -523 2262 -518
rect 2339 -526 2344 -521
rect 564 -548 569 -543
rect 443 -590 448 -585
rect 585 -605 590 -600
rect 806 -589 810 -584
rect 824 -589 828 -584
rect 806 -606 811 -601
rect 823 -606 828 -601
rect 962 -589 966 -584
rect 980 -589 984 -584
rect 962 -606 967 -601
rect 979 -606 984 -601
rect 1112 -589 1116 -584
rect 1130 -589 1134 -584
rect 1112 -606 1117 -601
rect 1129 -606 1134 -601
rect 1268 -589 1272 -584
rect 1286 -589 1290 -584
rect 1268 -606 1273 -601
rect 1285 -606 1290 -601
rect 1514 -579 1518 -574
rect 1539 -579 1543 -574
rect 1514 -596 1518 -591
rect 1539 -596 1543 -591
rect 1753 -578 1757 -573
rect 1777 -578 1781 -573
rect 1753 -595 1757 -590
rect 1777 -595 1781 -590
rect 1986 -578 1990 -573
rect 2010 -578 2014 -573
rect 1986 -595 1990 -590
rect 2010 -595 2014 -590
rect 2207 -578 2211 -573
rect 2231 -578 2235 -573
rect 2207 -595 2211 -590
rect 2231 -595 2235 -590
rect 2313 -581 2317 -576
rect 2313 -598 2317 -593
rect 564 -639 569 -634
rect 564 -649 569 -644
rect 564 -659 569 -654
<< metal1 >>
rect 1051 282 1054 295
rect 964 267 1008 270
rect 964 262 967 267
rect 984 262 987 267
rect 1005 266 1008 267
rect 1005 263 1029 266
rect 1005 262 1008 263
rect 950 259 963 262
rect 944 256 963 259
rect 1026 259 1029 263
rect 944 203 947 256
rect 974 244 977 256
rect 994 244 997 256
rect 974 241 1032 244
rect 1005 227 1008 241
rect 1040 244 1043 251
rect 1051 244 1054 277
rect 1085 274 1088 286
rect 1040 241 1054 244
rect 1085 244 1088 269
rect 1130 267 1174 270
rect 1130 266 1133 267
rect 1109 263 1133 266
rect 1109 259 1112 263
rect 1130 262 1133 263
rect 1151 262 1154 267
rect 1171 262 1174 267
rect 1175 259 1188 262
rect 1175 256 1198 259
rect 1095 244 1098 251
rect 1085 241 1098 244
rect 1040 227 1043 241
rect 950 221 963 227
rect 906 200 947 203
rect 906 142 909 200
rect 953 174 956 221
rect 1095 227 1098 241
rect 1141 244 1144 256
rect 1161 244 1164 256
rect 1106 241 1164 244
rect 1130 227 1133 241
rect 1175 221 1188 227
rect 1026 213 1029 219
rect 1025 210 1029 213
rect 1109 213 1112 219
rect 1109 210 1122 213
rect 969 206 972 209
rect 964 203 972 206
rect 964 160 967 203
rect 979 174 982 209
rect 989 200 992 209
rect 999 206 1002 209
rect 999 203 1017 206
rect 989 197 1009 200
rect 1006 177 1009 197
rect 979 171 997 174
rect 994 165 997 171
rect 987 162 1011 165
rect 940 157 967 160
rect 940 132 943 157
rect 781 129 943 132
rect 958 148 979 151
rect 781 123 784 129
rect 774 120 798 123
rect 745 106 766 109
rect 745 48 748 106
rect 781 87 784 112
rect 806 106 815 109
rect 812 87 815 106
rect 772 86 784 87
rect 772 84 800 86
rect 781 83 800 84
rect 756 78 759 81
rect 756 68 759 71
rect 783 66 786 83
rect 811 76 815 87
rect 805 73 815 76
rect 783 63 800 66
rect 767 48 772 52
rect 745 45 772 48
rect 755 13 758 45
rect 767 39 772 45
rect 776 37 779 57
rect 811 55 815 73
rect 805 52 815 55
rect 811 42 815 52
rect 808 39 871 42
rect 906 41 909 120
rect 958 90 961 148
rect 994 129 997 154
rect 1025 151 1028 210
rect 1043 203 1116 206
rect 1113 160 1116 203
rect 1119 174 1122 210
rect 1136 196 1139 209
rect 1146 185 1149 209
rect 1156 183 1159 209
rect 1166 200 1169 209
rect 1156 180 1171 183
rect 1182 174 1185 221
rect 1195 198 1198 256
rect 1369 227 1372 233
rect 1119 171 1185 174
rect 1193 177 1325 180
rect 1113 157 1128 160
rect 1125 151 1128 157
rect 1019 148 1028 151
rect 1025 141 1028 148
rect 1118 148 1142 151
rect 1025 129 1028 135
rect 985 128 997 129
rect 985 126 1013 128
rect 994 125 1013 126
rect 969 120 972 123
rect 969 110 972 113
rect 996 108 999 125
rect 1024 118 1028 129
rect 1018 115 1028 118
rect 996 105 1013 108
rect 980 90 985 94
rect 958 87 985 90
rect 925 54 928 82
rect 968 55 971 87
rect 980 81 985 87
rect 989 79 992 99
rect 1024 97 1028 115
rect 1018 94 1028 97
rect 1024 84 1028 94
rect 1089 134 1110 137
rect 1089 88 1092 134
rect 1125 115 1128 140
rect 1156 137 1159 171
rect 1193 167 1196 177
rect 1322 171 1325 177
rect 1315 168 1339 171
rect 1168 164 1196 167
rect 1286 154 1307 157
rect 1150 134 1159 137
rect 1156 115 1159 134
rect 1116 114 1128 115
rect 1116 112 1144 114
rect 1125 111 1144 112
rect 1100 106 1103 109
rect 1100 96 1103 99
rect 1127 94 1130 111
rect 1155 104 1159 115
rect 1149 101 1159 104
rect 1127 91 1144 94
rect 1021 81 1028 84
rect 1072 85 1092 88
rect 989 76 993 79
rect 990 69 993 76
rect 983 66 1007 69
rect 968 52 975 55
rect 968 41 971 52
rect 990 46 993 58
rect 1021 55 1024 81
rect 1015 52 1024 55
rect 776 34 780 37
rect 777 27 780 34
rect 770 24 794 27
rect 755 10 762 13
rect 755 3 758 10
rect 777 4 780 16
rect 808 13 811 39
rect 802 10 811 13
rect 755 0 762 3
rect 759 -3 762 0
rect 775 1 780 4
rect 775 -96 778 1
rect 808 -5 811 10
rect 837 -14 840 26
rect 830 -17 854 -14
rect 787 -31 822 -28
rect 801 -89 804 -31
rect 837 -50 840 -25
rect 868 -28 871 39
rect 862 -31 871 -28
rect 868 -50 871 -31
rect 828 -51 840 -50
rect 828 -53 856 -51
rect 837 -54 856 -53
rect 812 -59 815 -56
rect 812 -69 815 -66
rect 839 -71 842 -54
rect 867 -61 871 -50
rect 861 -64 871 -61
rect 839 -74 856 -71
rect 823 -89 828 -85
rect 791 -96 794 -90
rect 801 -92 828 -89
rect 775 -99 794 -96
rect 791 -144 794 -99
rect 811 -124 814 -92
rect 823 -98 828 -92
rect 832 -100 835 -80
rect 867 -82 871 -64
rect 889 38 971 41
rect 988 43 993 46
rect 889 -23 892 38
rect 925 -9 928 28
rect 956 24 980 27
rect 918 -12 942 -9
rect 889 -26 910 -23
rect 861 -85 871 -82
rect 889 -84 892 -26
rect 925 -45 928 -20
rect 956 -23 959 24
rect 950 -26 959 -23
rect 956 -45 959 -26
rect 916 -46 928 -45
rect 916 -48 944 -46
rect 925 -49 944 -48
rect 900 -54 903 -51
rect 900 -64 903 -61
rect 927 -66 930 -49
rect 955 -56 959 -45
rect 949 -59 959 -56
rect 927 -69 944 -66
rect 911 -84 916 -80
rect 867 -95 871 -85
rect 864 -98 871 -95
rect 832 -103 836 -100
rect 833 -110 836 -103
rect 826 -113 850 -110
rect 811 -127 818 -124
rect 811 -142 814 -127
rect 833 -133 836 -121
rect 864 -124 867 -98
rect 858 -127 867 -124
rect 831 -136 836 -133
rect 789 -147 794 -144
rect 789 -159 792 -147
rect 831 -151 834 -136
rect 800 -154 834 -151
rect 831 -157 834 -154
rect 789 -162 794 -159
rect 791 -224 794 -162
rect 735 -227 794 -224
rect 559 -247 715 -244
rect 559 -276 562 -247
rect 586 -253 647 -250
rect 586 -262 589 -253
rect 577 -265 605 -262
rect 550 -279 572 -276
rect 550 -295 553 -279
rect 586 -297 589 -273
rect 617 -276 620 -264
rect 610 -279 620 -276
rect 577 -298 589 -297
rect 577 -300 605 -298
rect 586 -301 605 -300
rect 539 -306 564 -303
rect 444 -316 564 -313
rect 444 -533 447 -316
rect 588 -318 591 -301
rect 617 -308 620 -279
rect 610 -311 620 -308
rect 588 -321 605 -318
rect 486 -326 564 -323
rect 486 -426 489 -326
rect 617 -329 620 -311
rect 610 -332 620 -329
rect 550 -341 553 -334
rect 572 -341 577 -332
rect 550 -344 577 -341
rect 558 -389 561 -344
rect 617 -347 620 -332
rect 644 -345 647 -253
rect 712 -337 715 -247
rect 657 -340 667 -337
rect 644 -348 650 -345
rect 644 -363 650 -362
rect 586 -365 650 -363
rect 586 -366 647 -365
rect 586 -375 589 -366
rect 577 -378 605 -375
rect 617 -379 620 -376
rect 657 -379 660 -340
rect 707 -340 715 -337
rect 691 -356 699 -353
rect 691 -369 694 -356
rect 675 -372 694 -369
rect 712 -369 715 -340
rect 707 -372 715 -369
rect 617 -383 660 -379
rect 550 -392 572 -389
rect 550 -408 553 -392
rect 586 -410 589 -386
rect 617 -389 620 -383
rect 610 -392 620 -389
rect 577 -411 589 -410
rect 577 -413 605 -411
rect 586 -414 605 -413
rect 513 -419 564 -416
rect 486 -429 564 -426
rect 486 -473 489 -429
rect 588 -431 591 -414
rect 617 -421 620 -392
rect 657 -395 660 -383
rect 657 -398 667 -395
rect 691 -401 694 -372
rect 712 -395 715 -372
rect 707 -398 715 -395
rect 675 -413 699 -410
rect 610 -424 620 -421
rect 588 -434 605 -431
rect 521 -439 564 -436
rect 455 -487 458 -473
rect 470 -476 498 -473
rect 455 -490 465 -487
rect 455 -496 458 -490
rect 444 -579 447 -538
rect 486 -543 489 -484
rect 503 -490 513 -487
rect 506 -497 509 -490
rect 505 -500 509 -497
rect 435 -582 463 -579
rect 425 -596 430 -593
rect 425 -605 428 -596
rect 444 -613 447 -590
rect 475 -593 478 -580
rect 468 -596 478 -593
rect 475 -603 478 -596
rect 444 -654 447 -618
rect 486 -644 489 -548
rect 505 -605 508 -500
rect 522 -579 525 -439
rect 617 -442 620 -424
rect 691 -422 694 -413
rect 691 -425 721 -422
rect 610 -445 620 -442
rect 550 -452 553 -447
rect 572 -452 577 -445
rect 550 -455 577 -452
rect 562 -497 565 -455
rect 617 -460 620 -445
rect 586 -474 706 -471
rect 586 -483 589 -474
rect 577 -486 605 -483
rect 550 -500 572 -497
rect 550 -503 553 -500
rect 586 -518 589 -494
rect 617 -497 620 -489
rect 610 -500 620 -497
rect 577 -519 589 -518
rect 577 -521 605 -519
rect 586 -522 605 -521
rect 539 -527 564 -524
rect 539 -537 564 -534
rect 588 -539 591 -522
rect 617 -529 620 -500
rect 610 -532 620 -529
rect 588 -542 605 -539
rect 539 -547 564 -544
rect 617 -550 620 -532
rect 610 -553 620 -550
rect 550 -558 553 -555
rect 572 -558 577 -553
rect 550 -561 577 -558
rect 558 -575 561 -561
rect 617 -567 620 -553
rect 703 -560 706 -474
rect 718 -550 721 -425
rect 735 -437 738 -227
rect 815 -237 818 -180
rect 864 -201 867 -127
rect 835 -204 867 -201
rect 835 -230 838 -204
rect 753 -240 818 -237
rect 753 -296 756 -240
rect 879 -247 882 -85
rect 889 -87 916 -84
rect 899 -119 902 -87
rect 911 -93 916 -87
rect 920 -95 923 -75
rect 955 -77 959 -59
rect 949 -80 959 -77
rect 955 -90 959 -80
rect 952 -93 959 -90
rect 920 -98 924 -95
rect 921 -105 924 -98
rect 914 -108 938 -105
rect 899 -122 906 -119
rect 899 -127 902 -122
rect 899 -130 903 -127
rect 921 -128 924 -116
rect 952 -119 955 -93
rect 946 -122 955 -119
rect 900 -133 903 -130
rect 919 -131 924 -128
rect 919 -145 922 -131
rect 952 -136 955 -122
rect 988 -170 991 43
rect 1021 27 1024 52
rect 1001 24 1024 27
rect 1072 -13 1075 85
rect 1089 76 1092 85
rect 1111 76 1116 80
rect 1079 19 1082 75
rect 1089 73 1116 76
rect 1099 41 1102 73
rect 1111 67 1116 73
rect 1120 65 1123 85
rect 1155 83 1159 101
rect 1149 80 1159 83
rect 1155 70 1159 80
rect 1152 67 1159 70
rect 1120 62 1124 65
rect 1121 55 1124 62
rect 1114 52 1138 55
rect 1099 38 1106 41
rect 1099 23 1102 38
rect 1121 32 1124 44
rect 1152 41 1155 67
rect 1188 47 1191 150
rect 1286 96 1289 154
rect 1322 135 1325 160
rect 1347 154 1356 157
rect 1353 135 1356 154
rect 1313 134 1325 135
rect 1313 132 1341 134
rect 1322 131 1341 132
rect 1297 126 1300 129
rect 1297 116 1300 119
rect 1324 114 1327 131
rect 1352 124 1356 135
rect 1346 121 1356 124
rect 1324 111 1341 114
rect 1308 96 1313 100
rect 1286 93 1313 96
rect 1296 61 1299 93
rect 1308 87 1313 93
rect 1317 85 1320 105
rect 1352 103 1356 121
rect 1346 100 1356 103
rect 1352 90 1356 100
rect 1349 87 1356 90
rect 1317 82 1321 85
rect 1318 75 1321 82
rect 1311 72 1335 75
rect 1296 58 1303 61
rect 1296 47 1299 58
rect 1318 52 1321 64
rect 1349 61 1352 87
rect 1343 58 1352 61
rect 1188 44 1299 47
rect 1316 49 1321 52
rect 1146 38 1155 41
rect 1119 29 1124 32
rect 1079 16 1113 19
rect 1110 -4 1113 16
rect 1119 6 1122 29
rect 1152 24 1155 38
rect 1152 23 1187 24
rect 1152 21 1183 23
rect 1172 12 1175 13
rect 1153 9 1175 12
rect 1153 0 1156 9
rect 1146 -3 1170 0
rect 1103 -7 1113 -4
rect 1092 -14 1095 -8
rect 1088 -17 1095 -14
rect 1088 -83 1091 -17
rect 1103 -27 1106 -7
rect 1114 -17 1138 -14
rect 1117 -22 1120 -17
rect 1116 -25 1120 -22
rect 1103 -30 1113 -27
rect 1101 -83 1104 -76
rect 1088 -86 1104 -83
rect 896 -173 991 -170
rect 988 -180 1034 -178
rect 1101 -180 1104 -86
rect 1110 -132 1113 -30
rect 1117 -75 1120 -25
rect 1153 -36 1156 -11
rect 1184 -14 1187 18
rect 1178 -17 1187 -14
rect 1233 -16 1236 44
rect 1254 35 1296 38
rect 1316 29 1319 49
rect 1349 46 1352 58
rect 1303 26 1319 29
rect 1322 43 1352 46
rect 1258 20 1261 23
rect 1255 17 1261 20
rect 1255 -2 1258 17
rect 1303 11 1306 26
rect 1322 23 1325 43
rect 1302 8 1306 11
rect 1248 -5 1272 -2
rect 1184 -36 1187 -17
rect 1144 -37 1156 -36
rect 1144 -39 1172 -37
rect 1153 -40 1172 -39
rect 1128 -45 1131 -42
rect 1128 -55 1131 -52
rect 1155 -57 1158 -40
rect 1183 -47 1187 -36
rect 1177 -50 1187 -47
rect 1155 -60 1172 -57
rect 1139 -75 1144 -71
rect 1117 -78 1144 -75
rect 1127 -110 1130 -78
rect 1139 -84 1144 -78
rect 1148 -86 1151 -66
rect 1183 -68 1187 -50
rect 1177 -71 1187 -68
rect 1183 -81 1187 -71
rect 1219 -19 1240 -16
rect 1219 -77 1222 -19
rect 1255 -38 1258 -13
rect 1280 -19 1289 -16
rect 1286 -38 1289 -19
rect 1246 -39 1258 -38
rect 1246 -41 1274 -39
rect 1255 -42 1274 -41
rect 1230 -47 1233 -44
rect 1230 -57 1233 -54
rect 1257 -59 1260 -42
rect 1285 -49 1289 -38
rect 1279 -52 1289 -49
rect 1257 -62 1274 -59
rect 1241 -77 1246 -73
rect 1180 -84 1187 -81
rect 1148 -89 1152 -86
rect 1149 -96 1152 -89
rect 1142 -99 1166 -96
rect 1127 -113 1134 -110
rect 1127 -124 1130 -113
rect 1149 -119 1152 -107
rect 1180 -110 1183 -84
rect 1174 -113 1183 -110
rect 1147 -122 1152 -119
rect 1147 -132 1150 -122
rect 1180 -126 1183 -113
rect 1110 -136 1150 -132
rect 1147 -139 1150 -136
rect 1127 -174 1130 -151
rect 988 -181 1104 -180
rect 988 -189 991 -181
rect 1031 -183 1104 -181
rect 1118 -177 1130 -174
rect 983 -192 1007 -189
rect 968 -207 975 -204
rect 775 -250 961 -247
rect 775 -281 778 -250
rect 768 -284 792 -281
rect 753 -299 760 -296
rect 753 -377 756 -299
rect 775 -342 778 -293
rect 800 -299 809 -296
rect 806 -309 809 -299
rect 835 -309 838 -260
rect 782 -312 845 -309
rect 782 -333 785 -312
rect 796 -318 799 -312
rect 828 -318 831 -312
rect 812 -342 815 -326
rect 775 -345 815 -342
rect 796 -350 799 -345
rect 832 -361 835 -358
rect 803 -369 806 -365
rect 745 -380 756 -377
rect 766 -372 806 -369
rect 820 -369 823 -365
rect 820 -372 859 -369
rect 745 -422 748 -380
rect 766 -383 769 -372
rect 856 -383 859 -372
rect 761 -386 777 -383
rect 758 -422 761 -418
rect 745 -425 761 -422
rect 758 -428 761 -425
rect 765 -431 769 -394
rect 774 -399 777 -386
rect 793 -386 802 -383
rect 799 -390 802 -386
rect 823 -386 832 -383
rect 799 -393 809 -390
rect 774 -402 785 -399
rect 799 -415 802 -393
rect 823 -390 826 -386
rect 848 -386 864 -383
rect 814 -393 826 -390
rect 793 -418 802 -415
rect 805 -414 809 -411
rect 816 -414 820 -411
rect 805 -417 820 -414
rect 823 -415 826 -393
rect 848 -399 851 -386
rect 840 -402 851 -399
rect 765 -434 781 -431
rect 778 -437 781 -434
rect 799 -437 802 -418
rect 811 -429 814 -417
rect 823 -418 832 -415
rect 855 -429 858 -394
rect 864 -423 867 -418
rect 811 -432 843 -429
rect 735 -440 781 -437
rect 778 -470 781 -440
rect 794 -440 829 -437
rect 794 -446 797 -440
rect 826 -446 829 -440
rect 810 -470 813 -454
rect 840 -470 843 -432
rect 778 -473 786 -470
rect 783 -497 786 -473
rect 810 -473 843 -470
rect 846 -432 858 -429
rect 846 -437 849 -432
rect 883 -437 886 -280
rect 846 -440 886 -437
rect 892 -437 895 -280
rect 900 -296 903 -262
rect 931 -267 961 -264
rect 931 -281 934 -267
rect 968 -272 971 -207
rect 988 -240 991 -201
rect 1015 -207 1024 -204
rect 1021 -220 1024 -207
rect 1021 -240 1024 -225
rect 983 -243 991 -240
rect 988 -256 991 -243
rect 1015 -243 1024 -240
rect 988 -259 1007 -256
rect 968 -275 975 -272
rect 1021 -272 1024 -243
rect 1031 -247 1034 -183
rect 1118 -204 1121 -177
rect 1209 -178 1212 -78
rect 1219 -80 1246 -77
rect 1138 -181 1212 -178
rect 1229 -112 1232 -80
rect 1241 -86 1246 -80
rect 1250 -88 1253 -68
rect 1285 -70 1289 -52
rect 1279 -73 1289 -70
rect 1285 -83 1289 -73
rect 1282 -86 1289 -83
rect 1250 -91 1254 -88
rect 1251 -98 1254 -91
rect 1244 -101 1268 -98
rect 1229 -115 1236 -112
rect 1138 -189 1141 -181
rect 1133 -192 1157 -189
rect 1118 -207 1125 -204
rect 1031 -250 1111 -247
rect 1081 -267 1111 -264
rect 1015 -275 1026 -272
rect 924 -284 948 -281
rect 968 -290 971 -275
rect 1023 -282 1026 -275
rect 1081 -281 1084 -267
rect 1118 -272 1121 -207
rect 1138 -240 1141 -201
rect 1165 -207 1174 -204
rect 1171 -240 1174 -207
rect 1133 -243 1141 -240
rect 1138 -256 1141 -243
rect 1165 -243 1174 -240
rect 1138 -259 1157 -256
rect 1118 -275 1125 -272
rect 1171 -272 1174 -243
rect 1177 -247 1180 -181
rect 1229 -204 1232 -115
rect 1251 -121 1254 -109
rect 1282 -112 1285 -86
rect 1276 -115 1285 -112
rect 1249 -124 1254 -121
rect 1249 -136 1252 -124
rect 1282 -156 1285 -115
rect 1302 -165 1305 8
rect 1322 -157 1325 18
rect 1316 -160 1325 -157
rect 1244 -168 1305 -165
rect 1285 -189 1288 -181
rect 1280 -192 1304 -189
rect 1322 -201 1325 -160
rect 1369 -172 1372 222
rect 1471 155 1474 427
rect 1478 359 1481 427
rect 1485 365 1488 427
rect 1492 372 1495 427
rect 1499 378 1502 427
rect 1499 375 2059 378
rect 1492 369 1929 372
rect 1485 362 1780 365
rect 1478 356 1649 359
rect 1543 349 1622 352
rect 1543 324 1546 349
rect 1550 344 1553 349
rect 1582 344 1585 349
rect 1608 344 1611 349
rect 1566 331 1569 336
rect 1566 328 1614 331
rect 1492 321 1546 324
rect 1455 152 1479 155
rect 1437 137 1447 140
rect 1437 130 1440 137
rect 1437 127 1463 130
rect 1418 104 1430 107
rect 1418 28 1421 104
rect 1424 87 1430 90
rect 1424 36 1427 87
rect 1437 82 1440 127
rect 1471 114 1474 143
rect 1492 140 1495 321
rect 1582 312 1585 328
rect 1623 331 1626 336
rect 1646 331 1649 356
rect 1684 349 1731 352
rect 1690 344 1693 349
rect 1710 344 1713 349
rect 1728 348 1731 349
rect 1745 348 1761 351
rect 1728 345 1748 348
rect 1675 338 1689 344
rect 1745 341 1748 345
rect 1623 328 1649 331
rect 1623 312 1626 328
rect 1700 326 1703 338
rect 1720 326 1723 338
rect 1700 323 1751 326
rect 1724 309 1727 323
rect 1759 326 1762 333
rect 1777 326 1780 362
rect 1834 351 1875 354
rect 1808 348 1816 351
rect 1813 346 1816 348
rect 1834 346 1837 351
rect 1854 346 1857 351
rect 1872 350 1875 351
rect 1872 347 1910 350
rect 1813 343 1833 346
rect 1819 340 1833 343
rect 1889 343 1892 347
rect 1759 323 1780 326
rect 1844 328 1847 340
rect 1864 328 1867 340
rect 1844 325 1895 328
rect 1759 309 1762 323
rect 1868 311 1871 325
rect 1903 328 1906 335
rect 1926 328 1929 369
rect 1977 352 2018 355
rect 1954 347 1966 350
rect 1977 347 1980 352
rect 1997 347 2000 352
rect 2015 351 2018 352
rect 2015 348 2035 351
rect 1962 341 1976 347
rect 2032 344 2035 348
rect 1903 325 1929 328
rect 1987 329 1990 341
rect 2007 329 2010 341
rect 1987 326 2038 329
rect 1903 311 1906 325
rect 2011 312 2014 326
rect 2046 329 2049 336
rect 2056 329 2059 375
rect 2046 326 2059 329
rect 2046 312 2049 326
rect 1550 297 1553 304
rect 1608 297 1611 304
rect 1675 303 1689 309
rect 1676 297 1679 303
rect 1550 294 1679 297
rect 1819 305 1833 311
rect 1558 265 1561 287
rect 1522 262 1561 265
rect 1522 172 1525 262
rect 1575 242 1578 287
rect 1550 205 1553 211
rect 1584 205 1587 294
rect 1676 285 1679 294
rect 1745 295 1748 301
rect 1736 292 1748 295
rect 1676 282 1682 285
rect 1695 269 1698 291
rect 1705 257 1708 291
rect 1715 265 1718 291
rect 1736 287 1739 292
rect 1820 287 1823 305
rect 1962 306 1976 312
rect 1889 297 1892 303
rect 1880 294 1892 297
rect 1736 285 1826 287
rect 1733 284 1826 285
rect 1733 282 1739 284
rect 1839 264 1842 293
rect 1705 254 1763 257
rect 1708 247 1727 250
rect 1529 202 1587 205
rect 1529 181 1532 202
rect 1543 196 1546 202
rect 1575 196 1578 202
rect 1559 172 1562 188
rect 1638 185 1712 188
rect 1638 182 1641 185
rect 1522 169 1562 172
rect 1543 164 1546 169
rect 1709 158 1712 185
rect 1760 175 1763 254
rect 1849 254 1852 293
rect 1859 264 1862 293
rect 1880 287 1883 294
rect 1963 288 1966 306
rect 2032 298 2035 304
rect 2023 295 2035 298
rect 1963 287 1969 288
rect 1877 285 1969 287
rect 1877 284 1966 285
rect 1982 278 1985 294
rect 1992 260 1995 294
rect 2002 279 2005 294
rect 2023 288 2026 295
rect 2020 285 2026 288
rect 1992 257 2234 260
rect 1849 250 1996 254
rect 1788 208 1791 211
rect 1767 205 1816 208
rect 1767 184 1770 205
rect 1781 199 1784 205
rect 1813 199 1816 205
rect 1797 175 1800 191
rect 1873 185 1945 188
rect 1873 182 1876 185
rect 1760 172 1800 175
rect 1781 167 1784 172
rect 1579 153 1582 156
rect 1693 155 1717 158
rect 1817 156 1820 159
rect 1942 158 1945 185
rect 1993 175 1996 250
rect 2021 208 2024 214
rect 2000 205 2049 208
rect 2000 184 2003 205
rect 2014 199 2017 205
rect 2046 199 2049 205
rect 2030 175 2033 191
rect 2109 188 2183 191
rect 2109 185 2112 188
rect 1993 172 2033 175
rect 2014 167 2017 172
rect 2180 161 2183 188
rect 2231 178 2234 257
rect 2259 211 2262 214
rect 2238 208 2287 211
rect 2238 187 2241 208
rect 2252 202 2255 208
rect 2284 202 2287 208
rect 2268 178 2271 194
rect 2231 175 2271 178
rect 2252 170 2255 175
rect 2367 170 2475 173
rect 1550 145 1553 149
rect 1487 137 1495 140
rect 1492 114 1495 137
rect 1513 142 1553 145
rect 1567 145 1570 149
rect 1788 148 1791 152
rect 1567 142 1606 145
rect 1513 131 1516 142
rect 1603 131 1606 142
rect 1675 140 1685 143
rect 1675 133 1678 140
rect 1508 128 1524 131
rect 1455 111 1474 114
rect 1471 98 1474 111
rect 1487 111 1495 114
rect 1471 95 1479 98
rect 1492 93 1495 111
rect 1505 93 1508 96
rect 1492 90 1508 93
rect 1437 79 1447 82
rect 1492 82 1495 90
rect 1505 87 1508 90
rect 1512 83 1516 120
rect 1521 115 1524 128
rect 1540 128 1549 131
rect 1546 124 1549 128
rect 1570 128 1579 131
rect 1546 121 1556 124
rect 1521 112 1532 115
rect 1546 99 1549 121
rect 1570 124 1573 128
rect 1595 128 1611 131
rect 1561 121 1573 124
rect 1540 96 1549 99
rect 1552 100 1556 103
rect 1563 100 1567 103
rect 1552 97 1567 100
rect 1570 99 1573 121
rect 1595 115 1598 128
rect 1675 130 1701 133
rect 1587 112 1598 115
rect 1487 79 1495 82
rect 1512 80 1528 83
rect 1437 57 1440 79
rect 1437 54 1454 57
rect 1451 51 1454 54
rect 1424 33 1461 36
rect 1418 25 1422 28
rect 1419 -105 1422 25
rect 1458 24 1461 33
rect 1442 21 1466 24
rect 1425 6 1434 9
rect 1425 -17 1428 6
rect 1451 -17 1454 -14
rect 1425 -20 1454 -17
rect 1425 -45 1428 -20
rect 1458 -45 1461 12
rect 1489 9 1492 79
rect 1525 44 1528 80
rect 1546 77 1549 96
rect 1558 85 1561 97
rect 1570 96 1579 99
rect 1602 85 1605 120
rect 1656 107 1668 110
rect 1611 91 1614 96
rect 1558 82 1590 85
rect 1541 74 1576 77
rect 1541 68 1544 74
rect 1573 68 1576 74
rect 1557 44 1560 60
rect 1587 44 1590 82
rect 1525 41 1533 44
rect 1530 17 1533 41
rect 1557 41 1590 44
rect 1593 82 1605 85
rect 1541 35 1544 38
rect 1573 35 1576 41
rect 1593 37 1596 82
rect 1579 34 1596 37
rect 1549 17 1552 20
rect 1530 14 1552 17
rect 1474 6 1492 9
rect 1425 -48 1434 -45
rect 1425 -77 1428 -48
rect 1458 -48 1466 -45
rect 1458 -61 1461 -48
rect 1442 -64 1461 -61
rect 1425 -80 1434 -77
rect 1478 -77 1481 6
rect 1549 -3 1552 14
rect 1503 -6 1552 -3
rect 1566 17 1569 20
rect 1579 17 1582 34
rect 1656 31 1659 107
rect 1662 90 1668 93
rect 1662 39 1665 90
rect 1675 85 1678 130
rect 1709 117 1712 146
rect 1751 145 1791 148
rect 1805 148 1808 152
rect 1926 155 1950 158
rect 2050 156 2053 159
rect 2164 158 2188 161
rect 2288 159 2291 162
rect 1805 145 1844 148
rect 2021 148 2024 152
rect 1725 140 1733 143
rect 1730 117 1733 140
rect 1751 134 1754 145
rect 1841 134 1844 145
rect 1908 140 1918 143
rect 1746 131 1762 134
rect 1693 114 1712 117
rect 1709 101 1712 114
rect 1725 114 1733 117
rect 1709 98 1717 101
rect 1730 96 1733 114
rect 1743 96 1746 99
rect 1730 93 1746 96
rect 1675 82 1685 85
rect 1730 85 1733 93
rect 1743 90 1746 93
rect 1750 86 1754 123
rect 1759 118 1762 131
rect 1778 131 1787 134
rect 1784 127 1787 131
rect 1808 131 1817 134
rect 1784 124 1794 127
rect 1759 115 1770 118
rect 1784 102 1787 124
rect 1808 127 1811 131
rect 1833 131 1849 134
rect 1799 124 1811 127
rect 1778 99 1787 102
rect 1790 103 1794 106
rect 1801 103 1805 106
rect 1790 100 1805 103
rect 1808 102 1811 124
rect 1833 118 1836 131
rect 1908 133 1911 140
rect 1908 130 1934 133
rect 1825 115 1836 118
rect 1725 82 1733 85
rect 1750 83 1766 86
rect 1675 60 1678 82
rect 1675 57 1692 60
rect 1689 54 1692 57
rect 1662 36 1699 39
rect 1656 28 1660 31
rect 1566 14 1582 17
rect 1488 -55 1495 -52
rect 1503 -64 1506 -6
rect 1566 -10 1569 14
rect 1522 -13 1569 -10
rect 1522 -52 1525 -13
rect 1529 -22 1578 -19
rect 1529 -43 1532 -22
rect 1543 -28 1546 -22
rect 1575 -28 1578 -22
rect 1559 -52 1562 -36
rect 1519 -55 1562 -52
rect 1492 -67 1506 -64
rect 1543 -60 1546 -55
rect 1492 -69 1495 -67
rect 1488 -72 1495 -69
rect 1579 -71 1582 -68
rect 1474 -80 1481 -77
rect 1478 -85 1481 -80
rect 1419 -108 1462 -105
rect 1459 -117 1462 -108
rect 1443 -120 1467 -117
rect 1492 -129 1495 -72
rect 1550 -79 1553 -75
rect 1513 -82 1553 -79
rect 1567 -79 1570 -75
rect 1567 -82 1606 -79
rect 1513 -93 1516 -82
rect 1603 -93 1606 -82
rect 1508 -96 1524 -93
rect 1426 -135 1435 -132
rect 1426 -147 1429 -135
rect 1426 -150 1442 -147
rect 1364 -175 1388 -172
rect 1349 -190 1356 -187
rect 1229 -207 1272 -204
rect 1177 -250 1258 -247
rect 1228 -267 1258 -264
rect 1165 -275 1176 -272
rect 1074 -284 1098 -281
rect 968 -293 1057 -290
rect 900 -299 916 -296
rect 909 -362 912 -299
rect 931 -342 934 -293
rect 1054 -296 1057 -293
rect 956 -299 965 -296
rect 1054 -299 1066 -296
rect 962 -309 965 -299
rect 938 -312 999 -309
rect 938 -333 941 -312
rect 952 -318 955 -312
rect 984 -318 987 -312
rect 968 -342 971 -326
rect 931 -345 971 -342
rect 952 -350 955 -345
rect 988 -361 991 -358
rect 903 -365 912 -362
rect 909 -377 912 -365
rect 959 -369 962 -365
rect 901 -380 912 -377
rect 922 -372 962 -369
rect 976 -369 979 -365
rect 976 -372 1015 -369
rect 901 -422 904 -380
rect 922 -383 925 -372
rect 1012 -383 1015 -372
rect 917 -386 933 -383
rect 914 -422 917 -418
rect 901 -425 917 -422
rect 914 -428 917 -425
rect 921 -431 925 -394
rect 930 -399 933 -386
rect 949 -386 958 -383
rect 955 -390 958 -386
rect 979 -386 988 -383
rect 955 -393 965 -390
rect 930 -402 941 -399
rect 955 -415 958 -393
rect 979 -390 982 -386
rect 1004 -386 1020 -383
rect 970 -393 982 -390
rect 949 -418 958 -415
rect 961 -414 965 -411
rect 972 -414 976 -411
rect 961 -417 976 -414
rect 979 -415 982 -393
rect 1004 -399 1007 -386
rect 996 -402 1007 -399
rect 921 -434 937 -431
rect 934 -437 937 -434
rect 955 -437 958 -418
rect 967 -429 970 -417
rect 979 -418 988 -415
rect 1011 -429 1014 -394
rect 1020 -423 1023 -418
rect 967 -432 999 -429
rect 892 -440 937 -437
rect 794 -479 797 -476
rect 826 -479 829 -473
rect 846 -477 849 -440
rect 934 -470 937 -440
rect 950 -440 985 -437
rect 950 -446 953 -440
rect 982 -446 985 -440
rect 966 -470 969 -454
rect 996 -470 999 -432
rect 934 -473 942 -470
rect 832 -480 849 -477
rect 802 -497 805 -494
rect 780 -500 805 -497
rect 819 -497 822 -494
rect 832 -497 835 -480
rect 939 -497 942 -473
rect 966 -473 999 -470
rect 1002 -432 1014 -429
rect 1002 -439 1005 -432
rect 1035 -439 1038 -304
rect 1002 -442 1038 -439
rect 1044 -437 1047 -304
rect 1059 -362 1062 -299
rect 1081 -342 1084 -293
rect 1118 -296 1121 -275
rect 1173 -282 1176 -275
rect 1228 -281 1231 -267
rect 1265 -272 1268 -207
rect 1285 -240 1288 -201
rect 1318 -204 1325 -201
rect 1312 -207 1321 -204
rect 1318 -240 1321 -207
rect 1332 -230 1335 -202
rect 1332 -233 1342 -230
rect 1280 -243 1288 -240
rect 1285 -256 1288 -243
rect 1312 -243 1321 -240
rect 1285 -259 1304 -256
rect 1265 -275 1272 -272
rect 1318 -272 1321 -243
rect 1312 -275 1321 -272
rect 1221 -284 1245 -281
rect 1106 -299 1115 -296
rect 1118 -299 1213 -296
rect 1112 -309 1115 -299
rect 1088 -312 1151 -309
rect 1088 -333 1091 -312
rect 1102 -318 1105 -312
rect 1134 -318 1137 -312
rect 1118 -342 1121 -326
rect 1081 -345 1121 -342
rect 1102 -350 1105 -345
rect 1138 -361 1141 -358
rect 1055 -365 1062 -362
rect 1059 -377 1062 -365
rect 1109 -369 1112 -365
rect 1051 -380 1062 -377
rect 1072 -372 1112 -369
rect 1126 -369 1129 -365
rect 1126 -372 1165 -369
rect 1051 -422 1054 -380
rect 1072 -383 1075 -372
rect 1162 -383 1165 -372
rect 1067 -386 1083 -383
rect 1064 -422 1067 -418
rect 1051 -425 1067 -422
rect 1064 -428 1067 -425
rect 1071 -431 1075 -394
rect 1080 -399 1083 -386
rect 1099 -386 1108 -383
rect 1105 -390 1108 -386
rect 1129 -386 1138 -383
rect 1105 -393 1115 -390
rect 1080 -402 1091 -399
rect 1105 -415 1108 -393
rect 1129 -390 1132 -386
rect 1154 -386 1170 -383
rect 1120 -393 1132 -390
rect 1099 -418 1108 -415
rect 1111 -414 1115 -411
rect 1122 -414 1126 -411
rect 1111 -417 1126 -414
rect 1129 -415 1132 -393
rect 1154 -399 1157 -386
rect 1146 -402 1157 -399
rect 1071 -434 1087 -431
rect 1084 -437 1087 -434
rect 1105 -437 1108 -418
rect 1117 -429 1120 -417
rect 1129 -418 1138 -415
rect 1161 -429 1164 -394
rect 1170 -423 1173 -418
rect 1117 -432 1149 -429
rect 1044 -440 1087 -437
rect 950 -479 953 -476
rect 982 -479 985 -473
rect 1002 -477 1005 -442
rect 1084 -470 1087 -440
rect 1100 -440 1135 -437
rect 1100 -446 1103 -440
rect 1132 -446 1135 -440
rect 1116 -470 1119 -454
rect 1146 -470 1149 -432
rect 1084 -473 1092 -470
rect 988 -480 1005 -477
rect 958 -497 961 -494
rect 819 -500 854 -497
rect 740 -527 743 -507
rect 780 -512 783 -500
rect 851 -512 854 -500
rect 936 -500 961 -497
rect 975 -497 978 -494
rect 988 -497 991 -480
rect 1089 -497 1092 -473
rect 1116 -473 1149 -470
rect 1152 -432 1164 -429
rect 1152 -437 1155 -432
rect 1183 -437 1186 -307
rect 1152 -440 1186 -437
rect 1192 -437 1195 -307
rect 1206 -362 1209 -299
rect 1228 -342 1231 -293
rect 1253 -299 1262 -296
rect 1259 -309 1262 -299
rect 1265 -297 1268 -275
rect 1265 -300 1271 -297
rect 1318 -309 1321 -275
rect 1331 -250 1342 -247
rect 1331 -275 1334 -250
rect 1349 -255 1352 -190
rect 1369 -223 1372 -184
rect 1402 -187 1405 -164
rect 1396 -190 1405 -187
rect 1402 -223 1405 -190
rect 1364 -226 1372 -223
rect 1369 -239 1372 -226
rect 1396 -226 1405 -223
rect 1369 -242 1388 -239
rect 1349 -258 1356 -255
rect 1402 -255 1405 -226
rect 1426 -186 1429 -150
rect 1459 -186 1462 -129
rect 1475 -135 1482 -132
rect 1479 -139 1482 -135
rect 1505 -139 1508 -128
rect 1479 -142 1508 -139
rect 1426 -189 1435 -186
rect 1426 -218 1429 -189
rect 1459 -189 1467 -186
rect 1459 -202 1462 -189
rect 1443 -205 1462 -202
rect 1426 -221 1435 -218
rect 1479 -218 1482 -142
rect 1505 -146 1508 -142
rect 1512 -141 1516 -104
rect 1521 -109 1524 -96
rect 1540 -96 1549 -93
rect 1546 -100 1549 -96
rect 1570 -96 1579 -93
rect 1546 -103 1556 -100
rect 1521 -112 1532 -109
rect 1546 -125 1549 -103
rect 1570 -100 1573 -96
rect 1595 -96 1611 -93
rect 1561 -103 1573 -100
rect 1540 -128 1549 -125
rect 1552 -124 1556 -121
rect 1563 -124 1567 -121
rect 1552 -127 1567 -124
rect 1570 -125 1573 -103
rect 1595 -109 1598 -96
rect 1587 -112 1598 -109
rect 1512 -144 1528 -141
rect 1525 -180 1528 -144
rect 1546 -147 1549 -128
rect 1558 -139 1561 -127
rect 1570 -128 1579 -125
rect 1602 -139 1605 -104
rect 1611 -133 1614 -128
rect 1558 -142 1590 -139
rect 1541 -150 1576 -147
rect 1541 -156 1544 -150
rect 1573 -156 1576 -150
rect 1557 -180 1560 -164
rect 1587 -180 1590 -142
rect 1525 -183 1533 -180
rect 1530 -193 1533 -183
rect 1557 -183 1590 -180
rect 1593 -142 1605 -139
rect 1489 -196 1533 -193
rect 1489 -213 1519 -210
rect 1530 -216 1533 -196
rect 1541 -189 1544 -186
rect 1573 -189 1576 -183
rect 1593 -187 1596 -142
rect 1579 -190 1596 -187
rect 1549 -216 1552 -204
rect 1566 -210 1569 -204
rect 1579 -210 1582 -190
rect 1562 -213 1582 -210
rect 1475 -221 1482 -218
rect 1426 -238 1429 -221
rect 1479 -226 1482 -221
rect 1530 -219 1552 -216
rect 1492 -236 1495 -223
rect 1396 -258 1405 -255
rect 1349 -261 1352 -258
rect 1402 -275 1405 -258
rect 1423 -241 1429 -238
rect 1458 -239 1495 -236
rect 1423 -275 1426 -241
rect 1458 -242 1461 -239
rect 1331 -278 1368 -275
rect 1402 -278 1426 -275
rect 1235 -312 1321 -309
rect 1235 -333 1238 -312
rect 1249 -318 1252 -312
rect 1281 -318 1284 -312
rect 1265 -342 1268 -326
rect 1228 -345 1268 -342
rect 1249 -350 1252 -345
rect 1285 -361 1288 -358
rect 1203 -365 1209 -362
rect 1206 -377 1209 -365
rect 1256 -369 1259 -365
rect 1198 -380 1209 -377
rect 1219 -372 1259 -369
rect 1273 -369 1276 -365
rect 1273 -372 1312 -369
rect 1198 -422 1201 -380
rect 1219 -383 1222 -372
rect 1309 -383 1312 -372
rect 1214 -386 1230 -383
rect 1211 -422 1214 -418
rect 1198 -425 1214 -422
rect 1211 -428 1214 -425
rect 1218 -431 1222 -394
rect 1227 -399 1230 -386
rect 1246 -386 1255 -383
rect 1252 -390 1255 -386
rect 1276 -386 1285 -383
rect 1252 -393 1262 -390
rect 1227 -402 1238 -399
rect 1252 -415 1255 -393
rect 1276 -390 1279 -386
rect 1301 -386 1317 -383
rect 1267 -393 1279 -390
rect 1246 -418 1255 -415
rect 1258 -414 1262 -411
rect 1269 -414 1273 -411
rect 1258 -417 1273 -414
rect 1276 -415 1279 -393
rect 1301 -399 1304 -386
rect 1293 -402 1304 -399
rect 1218 -434 1234 -431
rect 1231 -437 1234 -434
rect 1252 -437 1255 -418
rect 1264 -429 1267 -417
rect 1276 -418 1285 -415
rect 1308 -429 1311 -394
rect 1317 -423 1320 -418
rect 1264 -432 1296 -429
rect 1192 -440 1234 -437
rect 1100 -479 1103 -476
rect 1132 -479 1135 -473
rect 1152 -477 1155 -440
rect 1231 -470 1234 -440
rect 1247 -440 1282 -437
rect 1247 -446 1250 -440
rect 1279 -446 1282 -440
rect 1263 -470 1266 -454
rect 1293 -470 1296 -432
rect 1231 -473 1239 -470
rect 1138 -480 1155 -477
rect 1108 -497 1111 -494
rect 975 -500 1010 -497
rect 764 -515 788 -512
rect 846 -515 870 -512
rect 740 -530 756 -527
rect 653 -570 678 -567
rect 653 -575 656 -570
rect 558 -578 656 -575
rect 675 -575 678 -570
rect 675 -578 727 -575
rect 747 -578 750 -530
rect 780 -578 783 -524
rect 796 -530 804 -527
rect 831 -530 838 -527
rect 558 -608 561 -578
rect 664 -582 667 -578
rect 586 -585 667 -582
rect 586 -594 589 -585
rect 577 -597 605 -594
rect 550 -611 572 -608
rect 550 -625 553 -611
rect 586 -629 589 -605
rect 617 -608 620 -594
rect 610 -611 620 -608
rect 577 -630 589 -629
rect 577 -632 605 -630
rect 586 -633 605 -632
rect 538 -638 564 -635
rect 538 -648 564 -645
rect 444 -697 447 -659
rect 486 -690 489 -649
rect 588 -650 591 -633
rect 617 -640 620 -611
rect 723 -630 726 -578
rect 747 -581 756 -578
rect 747 -610 750 -581
rect 780 -581 788 -578
rect 780 -594 783 -581
rect 764 -597 783 -594
rect 747 -613 756 -610
rect 800 -610 803 -530
rect 810 -588 816 -585
rect 821 -588 824 -585
rect 796 -613 803 -610
rect 800 -630 803 -613
rect 807 -621 810 -606
rect 824 -621 827 -606
rect 831 -610 834 -530
rect 851 -578 854 -524
rect 894 -527 897 -507
rect 936 -512 939 -500
rect 1007 -512 1010 -500
rect 1086 -500 1111 -497
rect 1125 -497 1128 -494
rect 1138 -497 1141 -480
rect 1236 -497 1239 -473
rect 1263 -473 1296 -470
rect 1299 -432 1311 -429
rect 1299 -435 1302 -432
rect 1338 -435 1341 -293
rect 1299 -438 1341 -435
rect 1247 -479 1250 -476
rect 1279 -479 1282 -473
rect 1299 -477 1302 -438
rect 1285 -480 1302 -477
rect 1255 -497 1258 -494
rect 1125 -500 1160 -497
rect 1236 -500 1258 -497
rect 1272 -497 1275 -494
rect 1285 -497 1288 -480
rect 1272 -500 1316 -497
rect 920 -515 944 -512
rect 1002 -515 1026 -512
rect 878 -530 912 -527
rect 884 -578 887 -530
rect 846 -581 854 -578
rect 851 -594 854 -581
rect 878 -581 887 -578
rect 851 -597 870 -594
rect 831 -613 838 -610
rect 884 -610 887 -581
rect 878 -613 887 -610
rect 903 -578 906 -530
rect 936 -578 939 -524
rect 952 -530 960 -527
rect 987 -530 994 -527
rect 903 -581 912 -578
rect 903 -610 906 -581
rect 936 -581 944 -578
rect 936 -594 939 -581
rect 920 -597 939 -594
rect 903 -613 912 -610
rect 956 -610 959 -530
rect 966 -588 972 -585
rect 977 -588 980 -585
rect 952 -613 959 -610
rect 831 -630 834 -613
rect 956 -630 959 -613
rect 963 -621 966 -606
rect 980 -621 983 -606
rect 987 -610 990 -530
rect 1007 -578 1010 -524
rect 1047 -527 1050 -507
rect 1086 -512 1089 -500
rect 1157 -512 1160 -500
rect 1070 -515 1094 -512
rect 1152 -515 1176 -512
rect 1034 -530 1062 -527
rect 1040 -578 1043 -530
rect 1002 -581 1010 -578
rect 1007 -594 1010 -581
rect 1034 -581 1043 -578
rect 1007 -597 1026 -594
rect 987 -613 994 -610
rect 1040 -610 1043 -581
rect 1034 -613 1043 -610
rect 1053 -578 1056 -530
rect 1086 -578 1089 -524
rect 1102 -530 1110 -527
rect 1137 -530 1144 -527
rect 1053 -581 1062 -578
rect 1053 -610 1056 -581
rect 1086 -581 1094 -578
rect 1086 -594 1089 -581
rect 1070 -597 1089 -594
rect 1053 -613 1062 -610
rect 1106 -610 1109 -530
rect 1116 -588 1122 -585
rect 1127 -588 1130 -585
rect 1102 -613 1109 -610
rect 987 -630 990 -613
rect 1106 -630 1109 -613
rect 1113 -621 1116 -606
rect 1130 -621 1133 -606
rect 1137 -610 1140 -530
rect 1157 -578 1160 -524
rect 1199 -527 1202 -507
rect 1242 -512 1245 -500
rect 1313 -512 1316 -500
rect 1365 -510 1368 -278
rect 1423 -304 1426 -278
rect 1445 -245 1461 -242
rect 1445 -284 1448 -245
rect 1452 -254 1501 -251
rect 1452 -275 1455 -254
rect 1466 -260 1469 -254
rect 1498 -260 1501 -254
rect 1482 -284 1485 -268
rect 1445 -287 1485 -284
rect 1466 -292 1469 -287
rect 1502 -303 1505 -300
rect 1411 -307 1429 -304
rect 1411 -502 1414 -307
rect 1473 -311 1476 -307
rect 1436 -314 1476 -311
rect 1490 -311 1493 -307
rect 1490 -314 1529 -311
rect 1436 -325 1439 -314
rect 1526 -325 1529 -314
rect 1431 -328 1447 -325
rect 1428 -365 1431 -360
rect 1435 -373 1439 -336
rect 1444 -341 1447 -328
rect 1463 -328 1472 -325
rect 1469 -332 1472 -328
rect 1493 -328 1502 -325
rect 1469 -335 1479 -332
rect 1444 -344 1455 -341
rect 1469 -357 1472 -335
rect 1493 -332 1496 -328
rect 1518 -328 1534 -325
rect 1484 -335 1496 -332
rect 1463 -360 1472 -357
rect 1475 -356 1479 -353
rect 1486 -356 1490 -353
rect 1475 -359 1490 -356
rect 1493 -357 1496 -335
rect 1518 -341 1521 -328
rect 1510 -344 1521 -341
rect 1435 -376 1451 -373
rect 1448 -412 1451 -376
rect 1469 -379 1472 -360
rect 1481 -371 1484 -359
rect 1493 -360 1502 -357
rect 1525 -371 1528 -336
rect 1534 -365 1537 -360
rect 1481 -374 1513 -371
rect 1464 -382 1499 -379
rect 1464 -388 1467 -382
rect 1496 -388 1499 -382
rect 1480 -412 1483 -396
rect 1510 -412 1513 -374
rect 1448 -415 1456 -412
rect 1453 -439 1456 -415
rect 1480 -415 1513 -412
rect 1516 -374 1528 -371
rect 1464 -421 1467 -418
rect 1496 -421 1499 -415
rect 1516 -419 1519 -374
rect 1549 -406 1552 -219
rect 1502 -422 1519 -419
rect 1472 -439 1475 -436
rect 1453 -442 1475 -439
rect 1472 -458 1475 -442
rect 1489 -439 1492 -436
rect 1502 -439 1505 -422
rect 1489 -442 1505 -439
rect 1489 -493 1492 -442
rect 1488 -496 1492 -493
rect 1226 -515 1250 -512
rect 1308 -515 1332 -512
rect 1184 -530 1218 -527
rect 1190 -578 1193 -530
rect 1152 -581 1160 -578
rect 1157 -594 1160 -581
rect 1184 -581 1193 -578
rect 1157 -597 1176 -594
rect 1137 -613 1144 -610
rect 1190 -610 1193 -581
rect 1184 -613 1193 -610
rect 1209 -578 1212 -530
rect 1242 -578 1245 -524
rect 1258 -530 1266 -527
rect 1293 -530 1300 -527
rect 1209 -581 1218 -578
rect 1209 -610 1212 -581
rect 1242 -581 1250 -578
rect 1242 -594 1245 -581
rect 1226 -597 1245 -594
rect 1209 -613 1218 -610
rect 1262 -610 1265 -530
rect 1272 -588 1277 -585
rect 1282 -588 1286 -585
rect 1258 -613 1265 -610
rect 1137 -630 1140 -613
rect 1262 -630 1265 -613
rect 1269 -620 1272 -606
rect 1286 -620 1289 -606
rect 1293 -610 1296 -530
rect 1313 -578 1316 -524
rect 1411 -527 1414 -507
rect 1488 -512 1491 -496
rect 1566 -512 1569 -213
rect 1625 -235 1628 -87
rect 1657 -102 1660 28
rect 1696 27 1699 36
rect 1680 24 1704 27
rect 1663 9 1672 12
rect 1663 -14 1666 9
rect 1689 -14 1692 -11
rect 1663 -17 1692 -14
rect 1663 -42 1666 -17
rect 1696 -42 1699 15
rect 1727 12 1730 82
rect 1763 47 1766 83
rect 1784 80 1787 99
rect 1796 88 1799 100
rect 1808 99 1817 102
rect 1840 88 1843 123
rect 1889 107 1901 110
rect 1849 94 1852 99
rect 1796 85 1828 88
rect 1779 77 1814 80
rect 1779 71 1782 77
rect 1811 71 1814 77
rect 1795 47 1798 63
rect 1825 47 1828 85
rect 1763 44 1771 47
rect 1768 20 1771 44
rect 1795 44 1828 47
rect 1831 85 1843 88
rect 1779 38 1782 41
rect 1811 38 1814 44
rect 1831 40 1834 85
rect 1817 37 1834 40
rect 1787 20 1790 23
rect 1768 17 1790 20
rect 1712 9 1730 12
rect 1663 -45 1672 -42
rect 1663 -74 1666 -45
rect 1696 -45 1704 -42
rect 1696 -58 1699 -45
rect 1680 -61 1699 -58
rect 1663 -77 1672 -74
rect 1716 -74 1719 9
rect 1787 0 1790 17
rect 1741 -3 1790 0
rect 1804 20 1807 23
rect 1817 20 1820 37
rect 1889 31 1892 107
rect 1895 90 1901 93
rect 1895 39 1898 90
rect 1908 85 1911 130
rect 1942 117 1945 146
rect 1984 145 2024 148
rect 2038 148 2041 152
rect 2259 151 2262 155
rect 2038 145 2077 148
rect 1958 140 1966 143
rect 1963 117 1966 140
rect 1984 134 1987 145
rect 2074 134 2077 145
rect 2146 143 2156 146
rect 2146 136 2149 143
rect 1979 131 1995 134
rect 1926 114 1945 117
rect 1942 101 1945 114
rect 1958 114 1966 117
rect 1942 98 1950 101
rect 1963 96 1966 114
rect 1976 96 1979 99
rect 1963 93 1979 96
rect 1908 82 1918 85
rect 1963 85 1966 93
rect 1976 90 1979 93
rect 1983 86 1987 123
rect 1992 118 1995 131
rect 2011 131 2020 134
rect 2017 127 2020 131
rect 2041 131 2050 134
rect 2017 124 2027 127
rect 1992 115 2003 118
rect 2017 102 2020 124
rect 2041 127 2044 131
rect 2066 131 2082 134
rect 2032 124 2044 127
rect 2011 99 2020 102
rect 2023 103 2027 106
rect 2034 103 2038 106
rect 2023 100 2038 103
rect 2041 102 2044 124
rect 2066 118 2069 131
rect 2146 133 2172 136
rect 2058 115 2069 118
rect 1958 82 1966 85
rect 1983 83 1999 86
rect 1908 60 1911 82
rect 1908 57 1925 60
rect 1922 54 1925 57
rect 1895 36 1932 39
rect 1889 28 1893 31
rect 1804 17 1820 20
rect 1726 -52 1733 -49
rect 1741 -61 1744 -3
rect 1804 -7 1807 17
rect 1760 -10 1807 -7
rect 1760 -49 1763 -10
rect 1767 -19 1816 -16
rect 1767 -40 1770 -19
rect 1781 -25 1784 -19
rect 1813 -25 1816 -19
rect 1797 -49 1800 -33
rect 1757 -52 1800 -49
rect 1730 -64 1744 -61
rect 1781 -57 1784 -52
rect 1730 -66 1733 -64
rect 1726 -69 1733 -66
rect 1817 -68 1820 -65
rect 1712 -77 1719 -74
rect 1716 -82 1719 -77
rect 1657 -105 1700 -102
rect 1697 -114 1700 -105
rect 1681 -117 1705 -114
rect 1730 -126 1733 -69
rect 1788 -76 1791 -72
rect 1751 -79 1791 -76
rect 1805 -76 1808 -72
rect 1805 -79 1844 -76
rect 1751 -90 1754 -79
rect 1841 -90 1844 -79
rect 1746 -93 1762 -90
rect 1664 -132 1673 -129
rect 1664 -144 1667 -132
rect 1664 -147 1680 -144
rect 1664 -183 1667 -147
rect 1697 -183 1700 -126
rect 1713 -132 1720 -129
rect 1717 -136 1720 -132
rect 1743 -136 1746 -125
rect 1717 -139 1746 -136
rect 1664 -186 1673 -183
rect 1664 -215 1667 -186
rect 1697 -186 1705 -183
rect 1697 -199 1700 -186
rect 1681 -202 1700 -199
rect 1664 -218 1673 -215
rect 1717 -215 1720 -139
rect 1743 -143 1746 -139
rect 1750 -138 1754 -101
rect 1759 -106 1762 -93
rect 1778 -93 1787 -90
rect 1784 -97 1787 -93
rect 1808 -93 1817 -90
rect 1784 -100 1794 -97
rect 1759 -109 1770 -106
rect 1784 -122 1787 -100
rect 1808 -97 1811 -93
rect 1833 -93 1849 -90
rect 1799 -100 1811 -97
rect 1778 -125 1787 -122
rect 1790 -121 1794 -118
rect 1801 -121 1805 -118
rect 1790 -124 1805 -121
rect 1808 -122 1811 -100
rect 1833 -106 1836 -93
rect 1825 -109 1836 -106
rect 1750 -141 1766 -138
rect 1763 -177 1766 -141
rect 1784 -144 1787 -125
rect 1796 -136 1799 -124
rect 1808 -125 1817 -122
rect 1840 -136 1843 -101
rect 1849 -130 1852 -125
rect 1796 -139 1828 -136
rect 1779 -147 1814 -144
rect 1779 -153 1782 -147
rect 1811 -153 1814 -147
rect 1795 -177 1798 -161
rect 1825 -177 1828 -139
rect 1763 -180 1771 -177
rect 1768 -190 1771 -180
rect 1795 -180 1828 -177
rect 1831 -139 1843 -136
rect 1727 -193 1771 -190
rect 1727 -210 1757 -207
rect 1768 -213 1771 -193
rect 1779 -186 1782 -183
rect 1811 -186 1814 -180
rect 1831 -184 1834 -139
rect 1817 -187 1834 -184
rect 1787 -213 1790 -201
rect 1804 -207 1807 -201
rect 1817 -207 1820 -187
rect 1800 -210 1820 -207
rect 1713 -218 1720 -215
rect 1664 -235 1667 -218
rect 1717 -223 1720 -218
rect 1768 -216 1790 -213
rect 1730 -233 1733 -220
rect 1598 -238 1628 -235
rect 1661 -238 1667 -235
rect 1696 -236 1733 -233
rect 1598 -304 1601 -238
rect 1661 -301 1664 -238
rect 1696 -239 1699 -236
rect 1683 -242 1699 -239
rect 1683 -281 1686 -242
rect 1690 -251 1739 -248
rect 1690 -272 1693 -251
rect 1704 -257 1707 -251
rect 1736 -257 1739 -251
rect 1720 -281 1723 -265
rect 1683 -284 1723 -281
rect 1704 -289 1707 -284
rect 1740 -300 1743 -297
rect 1661 -304 1667 -301
rect 1595 -307 1601 -304
rect 1598 -360 1601 -307
rect 1711 -308 1714 -304
rect 1674 -311 1714 -308
rect 1728 -308 1731 -304
rect 1728 -311 1767 -308
rect 1674 -322 1677 -311
rect 1764 -322 1767 -311
rect 1669 -325 1685 -322
rect 1666 -360 1669 -357
rect 1598 -363 1669 -360
rect 1666 -366 1669 -363
rect 1673 -370 1677 -333
rect 1682 -338 1685 -325
rect 1701 -325 1710 -322
rect 1707 -329 1710 -325
rect 1731 -325 1740 -322
rect 1707 -332 1717 -329
rect 1682 -341 1693 -338
rect 1707 -354 1710 -332
rect 1731 -329 1734 -325
rect 1756 -325 1772 -322
rect 1722 -332 1734 -329
rect 1701 -357 1710 -354
rect 1713 -353 1717 -350
rect 1724 -353 1728 -350
rect 1713 -356 1728 -353
rect 1731 -354 1734 -332
rect 1756 -338 1759 -325
rect 1748 -341 1759 -338
rect 1673 -373 1689 -370
rect 1686 -409 1689 -373
rect 1707 -376 1710 -357
rect 1719 -368 1722 -356
rect 1731 -357 1740 -354
rect 1763 -368 1766 -333
rect 1772 -362 1775 -357
rect 1719 -371 1751 -368
rect 1702 -379 1737 -376
rect 1702 -385 1705 -379
rect 1734 -385 1737 -379
rect 1718 -409 1721 -393
rect 1748 -409 1751 -371
rect 1686 -412 1694 -409
rect 1691 -436 1694 -412
rect 1718 -412 1751 -409
rect 1754 -371 1766 -368
rect 1702 -418 1705 -415
rect 1734 -418 1737 -412
rect 1754 -416 1757 -371
rect 1787 -410 1790 -216
rect 1740 -419 1757 -416
rect 1710 -436 1713 -433
rect 1691 -439 1713 -436
rect 1710 -458 1713 -439
rect 1727 -436 1730 -433
rect 1740 -436 1743 -419
rect 1727 -439 1743 -436
rect 1472 -515 1496 -512
rect 1561 -515 1585 -512
rect 1340 -530 1464 -527
rect 1346 -578 1349 -530
rect 1365 -560 1368 -538
rect 1308 -581 1316 -578
rect 1313 -594 1316 -581
rect 1340 -581 1349 -578
rect 1313 -597 1332 -594
rect 1293 -613 1300 -610
rect 1346 -610 1349 -581
rect 1455 -568 1458 -530
rect 1488 -568 1491 -524
rect 1504 -530 1513 -527
rect 1540 -530 1553 -527
rect 1455 -571 1464 -568
rect 1455 -600 1458 -571
rect 1488 -571 1496 -568
rect 1488 -584 1491 -571
rect 1472 -587 1491 -584
rect 1455 -603 1464 -600
rect 1508 -600 1511 -530
rect 1518 -578 1526 -575
rect 1531 -578 1539 -575
rect 1518 -595 1524 -592
rect 1504 -603 1511 -600
rect 1521 -601 1524 -595
rect 1533 -595 1539 -592
rect 1533 -601 1536 -595
rect 1546 -600 1549 -530
rect 1566 -568 1569 -524
rect 1636 -527 1639 -506
rect 1727 -511 1730 -439
rect 1804 -511 1807 -210
rect 1863 -232 1866 -84
rect 1890 -102 1893 28
rect 1929 27 1932 36
rect 1913 24 1937 27
rect 1896 9 1905 12
rect 1896 -14 1899 9
rect 1922 -14 1925 -11
rect 1896 -17 1925 -14
rect 1896 -42 1899 -17
rect 1929 -42 1932 15
rect 1960 12 1963 82
rect 1996 47 1999 83
rect 2017 80 2020 99
rect 2029 88 2032 100
rect 2041 99 2050 102
rect 2073 88 2076 123
rect 2127 110 2139 113
rect 2082 94 2085 99
rect 2029 85 2061 88
rect 2012 77 2047 80
rect 2012 71 2015 77
rect 2044 71 2047 77
rect 2028 47 2031 63
rect 2058 47 2061 85
rect 1996 44 2004 47
rect 2001 20 2004 44
rect 2028 44 2061 47
rect 2064 85 2076 88
rect 2012 38 2015 41
rect 2044 38 2047 44
rect 2064 40 2067 85
rect 2050 37 2067 40
rect 2020 20 2023 23
rect 2001 17 2023 20
rect 1945 9 1963 12
rect 1896 -45 1905 -42
rect 1896 -74 1899 -45
rect 1929 -45 1937 -42
rect 1929 -58 1932 -45
rect 1913 -61 1932 -58
rect 1896 -77 1905 -74
rect 1949 -74 1952 9
rect 2020 0 2023 17
rect 1974 -3 2023 0
rect 2037 20 2040 23
rect 2050 20 2053 37
rect 2127 34 2130 110
rect 2133 93 2139 96
rect 2133 42 2136 93
rect 2146 88 2149 133
rect 2180 120 2183 149
rect 2222 148 2262 151
rect 2276 151 2279 155
rect 2276 148 2315 151
rect 2196 143 2204 146
rect 2201 120 2204 143
rect 2222 137 2225 148
rect 2312 137 2315 148
rect 2367 139 2370 170
rect 2400 154 2403 160
rect 2472 158 2475 170
rect 2461 155 2532 158
rect 2384 151 2408 154
rect 2461 149 2464 155
rect 2217 134 2233 137
rect 2164 117 2183 120
rect 2180 104 2183 117
rect 2196 117 2204 120
rect 2180 101 2188 104
rect 2201 99 2204 117
rect 2214 99 2217 102
rect 2201 96 2217 99
rect 2146 85 2156 88
rect 2201 88 2204 96
rect 2214 93 2217 96
rect 2221 89 2225 126
rect 2230 121 2233 134
rect 2249 134 2258 137
rect 2255 130 2258 134
rect 2279 134 2288 137
rect 2255 127 2265 130
rect 2230 118 2241 121
rect 2255 105 2258 127
rect 2279 130 2282 134
rect 2304 134 2320 137
rect 2270 127 2282 130
rect 2249 102 2258 105
rect 2261 106 2265 109
rect 2272 106 2276 109
rect 2261 103 2276 106
rect 2279 105 2282 127
rect 2304 121 2307 134
rect 2367 136 2376 139
rect 2296 118 2307 121
rect 2196 85 2204 88
rect 2221 86 2237 89
rect 2146 63 2149 85
rect 2146 60 2163 63
rect 2160 57 2163 60
rect 2133 39 2170 42
rect 2127 31 2131 34
rect 2037 17 2053 20
rect 1959 -52 1966 -49
rect 1974 -61 1977 -3
rect 2037 -7 2040 17
rect 1993 -10 2040 -7
rect 1993 -49 1996 -10
rect 2000 -19 2049 -16
rect 2000 -40 2003 -19
rect 2014 -25 2017 -19
rect 2046 -25 2049 -19
rect 2030 -49 2033 -33
rect 1990 -52 2033 -49
rect 1963 -64 1977 -61
rect 2014 -57 2017 -52
rect 1963 -66 1966 -64
rect 1959 -69 1966 -66
rect 2050 -68 2053 -65
rect 1945 -77 1952 -74
rect 1949 -82 1952 -77
rect 1890 -105 1933 -102
rect 1930 -114 1933 -105
rect 1914 -117 1938 -114
rect 1963 -126 1966 -69
rect 2021 -76 2024 -72
rect 1984 -79 2024 -76
rect 2038 -76 2041 -72
rect 2038 -79 2077 -76
rect 1984 -90 1987 -79
rect 2074 -90 2077 -79
rect 1979 -93 1995 -90
rect 1836 -235 1866 -232
rect 1897 -132 1906 -129
rect 1897 -144 1900 -132
rect 1897 -147 1913 -144
rect 1897 -183 1900 -147
rect 1930 -183 1933 -126
rect 1946 -132 1953 -129
rect 1950 -136 1953 -132
rect 1976 -136 1979 -125
rect 1950 -139 1979 -136
rect 1897 -186 1906 -183
rect 1897 -215 1900 -186
rect 1930 -186 1938 -183
rect 1930 -199 1933 -186
rect 1914 -202 1933 -199
rect 1897 -218 1906 -215
rect 1950 -215 1953 -139
rect 1976 -143 1979 -139
rect 1983 -138 1987 -101
rect 1992 -106 1995 -93
rect 2011 -93 2020 -90
rect 2017 -97 2020 -93
rect 2041 -93 2050 -90
rect 2017 -100 2027 -97
rect 1992 -109 2003 -106
rect 2017 -122 2020 -100
rect 2041 -97 2044 -93
rect 2066 -93 2082 -90
rect 2032 -100 2044 -97
rect 2011 -125 2020 -122
rect 2023 -121 2027 -118
rect 2034 -121 2038 -118
rect 2023 -124 2038 -121
rect 2041 -122 2044 -100
rect 2066 -106 2069 -93
rect 2058 -109 2069 -106
rect 1983 -141 1999 -138
rect 1996 -177 1999 -141
rect 2017 -144 2020 -125
rect 2029 -136 2032 -124
rect 2041 -125 2050 -122
rect 2073 -136 2076 -101
rect 2082 -130 2085 -125
rect 2029 -139 2061 -136
rect 2012 -147 2047 -144
rect 2012 -153 2015 -147
rect 2044 -153 2047 -147
rect 2028 -177 2031 -161
rect 2058 -177 2061 -139
rect 1996 -180 2004 -177
rect 2001 -190 2004 -180
rect 2028 -180 2061 -177
rect 2064 -139 2076 -136
rect 1960 -193 2004 -190
rect 1960 -210 1990 -207
rect 2001 -213 2004 -193
rect 2012 -186 2015 -183
rect 2044 -186 2047 -180
rect 2064 -184 2067 -139
rect 2050 -187 2067 -184
rect 2020 -213 2023 -201
rect 2037 -207 2040 -201
rect 2050 -207 2053 -187
rect 2033 -210 2053 -207
rect 1946 -218 1953 -215
rect 1897 -235 1900 -218
rect 1950 -223 1953 -218
rect 2001 -216 2023 -213
rect 1963 -233 1966 -220
rect 1836 -301 1839 -235
rect 1833 -304 1839 -301
rect 1894 -238 1900 -235
rect 1929 -236 1966 -233
rect 1894 -301 1897 -238
rect 1929 -239 1932 -236
rect 1916 -242 1932 -239
rect 1916 -281 1919 -242
rect 1923 -251 1972 -248
rect 1923 -272 1926 -251
rect 1937 -257 1940 -251
rect 1969 -257 1972 -251
rect 1953 -281 1956 -265
rect 1916 -284 1956 -281
rect 1937 -289 1940 -284
rect 1973 -300 1976 -297
rect 1894 -304 1900 -301
rect 1836 -361 1839 -304
rect 1944 -308 1947 -304
rect 1907 -311 1947 -308
rect 1961 -308 1964 -304
rect 1961 -311 2000 -308
rect 1907 -322 1910 -311
rect 1997 -322 2000 -311
rect 1902 -325 1918 -322
rect 1899 -361 1902 -357
rect 1836 -364 1902 -361
rect 1836 -365 1839 -364
rect 1899 -367 1902 -364
rect 1906 -370 1910 -333
rect 1915 -338 1918 -325
rect 1934 -325 1943 -322
rect 1940 -329 1943 -325
rect 1964 -325 1973 -322
rect 1940 -332 1950 -329
rect 1915 -341 1926 -338
rect 1940 -354 1943 -332
rect 1964 -329 1967 -325
rect 1989 -325 2005 -322
rect 1955 -332 1967 -329
rect 1934 -357 1943 -354
rect 1946 -353 1950 -350
rect 1957 -353 1961 -350
rect 1946 -356 1961 -353
rect 1964 -354 1967 -332
rect 1989 -338 1992 -325
rect 1981 -341 1992 -338
rect 1906 -373 1922 -370
rect 1919 -409 1922 -373
rect 1940 -376 1943 -357
rect 1952 -368 1955 -356
rect 1964 -357 1973 -354
rect 1996 -368 1999 -333
rect 2005 -362 2008 -357
rect 1952 -371 1984 -368
rect 1935 -379 1970 -376
rect 1935 -385 1938 -379
rect 1967 -385 1970 -379
rect 1951 -409 1954 -393
rect 1981 -409 1984 -371
rect 1919 -412 1927 -409
rect 1924 -436 1927 -412
rect 1951 -412 1984 -409
rect 1987 -371 1999 -368
rect 1935 -418 1938 -415
rect 1967 -418 1970 -412
rect 1987 -416 1990 -371
rect 2020 -409 2023 -216
rect 1973 -419 1990 -416
rect 1943 -436 1946 -433
rect 1924 -439 1946 -436
rect 1943 -458 1946 -439
rect 1960 -436 1963 -433
rect 1973 -436 1976 -419
rect 1960 -439 1976 -436
rect 1711 -514 1735 -511
rect 1799 -514 1823 -511
rect 1694 -527 1703 -526
rect 1593 -529 1703 -527
rect 1593 -530 1697 -529
rect 1599 -568 1602 -530
rect 1561 -571 1569 -568
rect 1566 -584 1569 -571
rect 1593 -571 1602 -568
rect 1566 -587 1585 -584
rect 1340 -613 1349 -610
rect 1293 -630 1296 -613
rect 1508 -614 1511 -603
rect 1546 -603 1553 -600
rect 1599 -600 1602 -571
rect 1593 -603 1602 -600
rect 1694 -567 1697 -530
rect 1727 -567 1730 -523
rect 1743 -529 1754 -526
rect 1781 -529 1791 -526
rect 1694 -570 1703 -567
rect 1694 -599 1697 -570
rect 1727 -570 1735 -567
rect 1727 -583 1730 -570
rect 1711 -586 1730 -583
rect 1694 -602 1703 -599
rect 1747 -599 1750 -529
rect 1757 -577 1765 -574
rect 1770 -577 1777 -574
rect 1757 -594 1763 -591
rect 1743 -602 1750 -599
rect 1760 -600 1763 -594
rect 1771 -594 1777 -591
rect 1771 -600 1774 -594
rect 1784 -599 1787 -529
rect 1804 -567 1807 -523
rect 1862 -526 1865 -506
rect 1960 -511 1963 -439
rect 2037 -511 2040 -210
rect 2096 -232 2099 -84
rect 2128 -99 2131 31
rect 2167 30 2170 39
rect 2151 27 2175 30
rect 2134 12 2143 15
rect 2134 -11 2137 12
rect 2160 -11 2163 -8
rect 2134 -14 2163 -11
rect 2134 -39 2137 -14
rect 2167 -39 2170 18
rect 2198 15 2201 85
rect 2234 50 2237 86
rect 2255 83 2258 102
rect 2267 91 2270 103
rect 2279 102 2288 105
rect 2311 91 2314 126
rect 2367 103 2370 136
rect 2400 103 2403 142
rect 2497 149 2500 155
rect 2529 149 2532 155
rect 2416 136 2423 139
rect 2320 97 2323 102
rect 2367 100 2376 103
rect 2267 88 2299 91
rect 2250 80 2285 83
rect 2250 74 2253 80
rect 2282 74 2285 80
rect 2266 50 2269 66
rect 2296 50 2299 88
rect 2234 47 2242 50
rect 2239 23 2242 47
rect 2266 47 2299 50
rect 2302 88 2314 91
rect 2250 41 2253 44
rect 2282 41 2285 47
rect 2302 43 2305 88
rect 2288 40 2305 43
rect 2367 71 2370 100
rect 2400 100 2408 103
rect 2400 87 2403 100
rect 2384 84 2403 87
rect 2420 88 2423 136
rect 2446 125 2449 141
rect 2434 122 2449 125
rect 2434 96 2437 122
rect 2446 117 2449 122
rect 2513 125 2516 141
rect 2458 122 2516 125
rect 2497 117 2500 122
rect 2430 93 2437 96
rect 2461 105 2464 109
rect 2529 105 2532 109
rect 2461 102 2545 105
rect 2461 88 2464 102
rect 2504 88 2507 95
rect 2521 91 2524 95
rect 2521 88 2530 91
rect 2420 85 2464 88
rect 2367 68 2376 71
rect 2420 71 2423 85
rect 2430 76 2437 79
rect 2416 68 2423 71
rect 2258 23 2261 26
rect 2239 20 2261 23
rect 2183 12 2201 15
rect 2134 -42 2143 -39
rect 2134 -71 2137 -42
rect 2167 -42 2175 -39
rect 2167 -55 2170 -42
rect 2151 -58 2170 -55
rect 2134 -74 2143 -71
rect 2187 -71 2190 12
rect 2258 3 2261 20
rect 2212 0 2261 3
rect 2275 23 2278 26
rect 2288 23 2291 40
rect 2275 20 2291 23
rect 2367 35 2370 68
rect 2420 63 2423 68
rect 2434 48 2437 76
rect 2504 75 2507 83
rect 2521 79 2530 82
rect 2521 75 2524 79
rect 2542 68 2545 102
rect 2461 65 2545 68
rect 2461 61 2464 65
rect 2529 61 2532 65
rect 2446 48 2449 53
rect 2434 45 2449 48
rect 2367 32 2431 35
rect 2197 -49 2204 -46
rect 2212 -58 2215 0
rect 2275 -4 2278 20
rect 2231 -7 2278 -4
rect 2231 -46 2234 -7
rect 2238 -16 2287 -13
rect 2238 -37 2241 -16
rect 2252 -22 2255 -16
rect 2284 -22 2287 -16
rect 2367 -20 2370 32
rect 2428 9 2431 32
rect 2446 29 2449 45
rect 2497 48 2500 53
rect 2458 45 2516 48
rect 2513 29 2516 45
rect 2461 15 2464 21
rect 2497 15 2500 21
rect 2529 15 2532 21
rect 2461 12 2532 15
rect 2461 9 2464 12
rect 2400 -5 2403 7
rect 2428 6 2464 9
rect 2461 -1 2464 6
rect 2461 -4 2532 -1
rect 2384 -8 2408 -5
rect 2461 -10 2464 -4
rect 2367 -23 2376 -20
rect 2268 -46 2271 -30
rect 2228 -49 2271 -46
rect 2201 -61 2215 -58
rect 2252 -54 2255 -49
rect 2201 -63 2204 -61
rect 2197 -66 2204 -63
rect 2288 -65 2291 -62
rect 2367 -56 2370 -23
rect 2400 -56 2403 -17
rect 2497 -10 2500 -4
rect 2529 -10 2532 -4
rect 2416 -23 2423 -20
rect 2367 -59 2376 -56
rect 2183 -74 2190 -71
rect 2187 -79 2190 -74
rect 2128 -102 2171 -99
rect 2168 -111 2171 -102
rect 2152 -114 2176 -111
rect 2201 -123 2204 -66
rect 2259 -73 2262 -69
rect 2222 -76 2262 -73
rect 2276 -73 2279 -69
rect 2276 -76 2315 -73
rect 2222 -87 2225 -76
rect 2312 -87 2315 -76
rect 2217 -90 2233 -87
rect 2135 -129 2144 -126
rect 2135 -141 2138 -129
rect 2135 -144 2151 -141
rect 2135 -180 2138 -144
rect 2168 -180 2171 -123
rect 2184 -129 2191 -126
rect 2188 -133 2191 -129
rect 2214 -133 2217 -122
rect 2188 -136 2217 -133
rect 2135 -183 2144 -180
rect 2135 -212 2138 -183
rect 2168 -183 2176 -180
rect 2168 -196 2171 -183
rect 2152 -199 2171 -196
rect 2135 -215 2144 -212
rect 2188 -212 2191 -136
rect 2214 -140 2217 -136
rect 2221 -135 2225 -98
rect 2230 -103 2233 -90
rect 2249 -90 2258 -87
rect 2255 -94 2258 -90
rect 2279 -90 2288 -87
rect 2255 -97 2265 -94
rect 2230 -106 2241 -103
rect 2255 -119 2258 -97
rect 2279 -94 2282 -90
rect 2304 -90 2320 -87
rect 2270 -97 2282 -94
rect 2249 -122 2258 -119
rect 2261 -118 2265 -115
rect 2272 -118 2276 -115
rect 2261 -121 2276 -118
rect 2279 -119 2282 -97
rect 2304 -103 2307 -90
rect 2296 -106 2307 -103
rect 2221 -138 2237 -135
rect 2234 -174 2237 -138
rect 2255 -141 2258 -122
rect 2267 -133 2270 -121
rect 2279 -122 2288 -119
rect 2311 -133 2314 -98
rect 2320 -127 2323 -122
rect 2267 -136 2299 -133
rect 2250 -144 2285 -141
rect 2250 -150 2253 -144
rect 2282 -150 2285 -144
rect 2266 -174 2269 -158
rect 2296 -174 2299 -136
rect 2234 -177 2242 -174
rect 2239 -187 2242 -177
rect 2266 -177 2299 -174
rect 2302 -136 2314 -133
rect 2198 -190 2242 -187
rect 2198 -207 2228 -204
rect 2239 -210 2242 -190
rect 2250 -183 2253 -180
rect 2282 -183 2285 -177
rect 2302 -181 2305 -136
rect 2288 -184 2305 -181
rect 2258 -210 2261 -198
rect 2275 -204 2278 -198
rect 2288 -204 2291 -184
rect 2271 -207 2291 -204
rect 2184 -215 2191 -212
rect 2135 -232 2138 -215
rect 2188 -220 2191 -215
rect 2239 -213 2261 -210
rect 2201 -230 2204 -217
rect 2069 -235 2099 -232
rect 2132 -235 2138 -232
rect 2167 -233 2204 -230
rect 2069 -301 2072 -235
rect 2132 -298 2135 -235
rect 2167 -236 2170 -233
rect 2154 -239 2170 -236
rect 2154 -278 2157 -239
rect 2161 -248 2210 -245
rect 2161 -269 2164 -248
rect 2175 -254 2178 -248
rect 2207 -254 2210 -248
rect 2191 -278 2194 -262
rect 2154 -281 2194 -278
rect 2175 -286 2178 -281
rect 2211 -297 2214 -294
rect 2132 -301 2138 -298
rect 2066 -304 2072 -301
rect 2069 -357 2072 -304
rect 2182 -305 2185 -301
rect 2145 -308 2185 -305
rect 2199 -305 2202 -301
rect 2199 -308 2238 -305
rect 2145 -319 2148 -308
rect 2235 -319 2238 -308
rect 2140 -322 2156 -319
rect 2137 -357 2140 -354
rect 2069 -360 2140 -357
rect 2137 -363 2140 -360
rect 2144 -367 2148 -330
rect 2153 -335 2156 -322
rect 2172 -322 2181 -319
rect 2178 -326 2181 -322
rect 2202 -322 2211 -319
rect 2178 -329 2188 -326
rect 2153 -338 2164 -335
rect 2178 -351 2181 -329
rect 2202 -326 2205 -322
rect 2227 -322 2243 -319
rect 2193 -329 2205 -326
rect 2172 -354 2181 -351
rect 2184 -350 2188 -347
rect 2195 -350 2199 -347
rect 2184 -353 2199 -350
rect 2202 -351 2205 -329
rect 2227 -335 2230 -322
rect 2219 -338 2230 -335
rect 2144 -370 2160 -367
rect 2157 -406 2160 -370
rect 2178 -373 2181 -354
rect 2190 -365 2193 -353
rect 2202 -354 2211 -351
rect 2234 -365 2237 -330
rect 2243 -359 2246 -354
rect 2190 -368 2222 -365
rect 2173 -376 2208 -373
rect 2173 -382 2176 -376
rect 2205 -382 2208 -376
rect 2189 -406 2192 -390
rect 2219 -406 2222 -368
rect 2157 -409 2165 -406
rect 2162 -433 2165 -409
rect 2189 -409 2222 -406
rect 2225 -368 2237 -365
rect 2173 -415 2176 -412
rect 2205 -415 2208 -409
rect 2225 -413 2228 -368
rect 2211 -416 2228 -413
rect 2181 -433 2184 -430
rect 2162 -436 2184 -433
rect 1944 -514 1968 -511
rect 2032 -514 2056 -511
rect 1831 -529 1936 -526
rect 1837 -567 1840 -529
rect 1799 -570 1807 -567
rect 1804 -583 1807 -570
rect 1831 -570 1840 -567
rect 1804 -586 1823 -583
rect 1546 -614 1549 -603
rect 1747 -614 1750 -602
rect 1784 -602 1791 -599
rect 1837 -599 1840 -570
rect 1831 -602 1840 -599
rect 1927 -567 1930 -529
rect 1960 -567 1963 -523
rect 1976 -529 1987 -526
rect 2014 -529 2024 -526
rect 1927 -570 1936 -567
rect 1927 -599 1930 -570
rect 1960 -570 1968 -567
rect 1960 -583 1963 -570
rect 1944 -586 1963 -583
rect 1927 -602 1936 -599
rect 1980 -599 1983 -529
rect 1990 -577 1998 -574
rect 2003 -577 2010 -574
rect 1990 -594 1996 -591
rect 1976 -602 1983 -599
rect 1993 -600 1996 -594
rect 2004 -594 2010 -591
rect 2004 -600 2007 -594
rect 2017 -599 2020 -529
rect 2037 -567 2040 -523
rect 2105 -526 2108 -506
rect 2181 -511 2184 -436
rect 2198 -433 2201 -430
rect 2211 -433 2214 -416
rect 2198 -436 2214 -433
rect 2198 -450 2201 -436
rect 2258 -511 2261 -213
rect 2275 -459 2278 -207
rect 2334 -229 2337 -81
rect 2367 -88 2370 -59
rect 2400 -59 2408 -56
rect 2400 -72 2403 -59
rect 2384 -75 2403 -72
rect 2420 -71 2423 -23
rect 2446 -34 2449 -18
rect 2434 -37 2449 -34
rect 2434 -63 2437 -37
rect 2446 -42 2449 -37
rect 2513 -34 2516 -18
rect 2542 -28 2545 65
rect 2458 -37 2516 -34
rect 2541 -31 2545 -28
rect 2497 -42 2500 -37
rect 2430 -66 2437 -63
rect 2461 -54 2464 -50
rect 2529 -54 2532 -50
rect 2541 -54 2544 -31
rect 2461 -57 2544 -54
rect 2461 -71 2464 -57
rect 2504 -70 2507 -64
rect 2521 -68 2524 -64
rect 2420 -74 2464 -71
rect 2307 -232 2337 -229
rect 2366 -91 2376 -88
rect 2420 -88 2423 -74
rect 2521 -71 2530 -68
rect 2430 -83 2437 -80
rect 2416 -91 2423 -88
rect 2366 -117 2369 -91
rect 2420 -96 2423 -91
rect 2434 -111 2437 -83
rect 2504 -84 2507 -75
rect 2521 -80 2530 -77
rect 2521 -84 2524 -80
rect 2541 -91 2544 -57
rect 2461 -94 2544 -91
rect 2461 -98 2464 -94
rect 2529 -98 2532 -94
rect 2446 -111 2449 -106
rect 2434 -114 2449 -111
rect 2366 -120 2432 -117
rect 2366 -174 2369 -120
rect 2429 -147 2432 -120
rect 2446 -130 2449 -114
rect 2497 -111 2500 -106
rect 2458 -114 2516 -111
rect 2513 -130 2516 -114
rect 2461 -144 2464 -138
rect 2497 -144 2500 -138
rect 2529 -144 2532 -138
rect 2461 -147 2532 -144
rect 2399 -159 2402 -147
rect 2429 -150 2465 -147
rect 2462 -155 2465 -150
rect 2460 -158 2531 -155
rect 2383 -162 2407 -159
rect 2460 -164 2463 -158
rect 2366 -177 2375 -174
rect 2366 -210 2369 -177
rect 2399 -210 2402 -171
rect 2496 -164 2499 -158
rect 2528 -164 2531 -158
rect 2415 -177 2422 -174
rect 2366 -213 2375 -210
rect 2307 -298 2310 -232
rect 2304 -301 2310 -298
rect 2307 -447 2310 -301
rect 2366 -242 2369 -213
rect 2399 -213 2407 -210
rect 2399 -226 2402 -213
rect 2383 -229 2402 -226
rect 2419 -226 2422 -177
rect 2445 -188 2448 -172
rect 2433 -191 2448 -188
rect 2433 -217 2436 -191
rect 2445 -196 2448 -191
rect 2512 -188 2515 -172
rect 2457 -191 2515 -188
rect 2496 -196 2499 -191
rect 2429 -220 2436 -217
rect 2460 -208 2463 -204
rect 2528 -208 2531 -204
rect 2541 -208 2544 -94
rect 2460 -211 2544 -208
rect 2460 -226 2463 -211
rect 2503 -225 2506 -218
rect 2520 -222 2523 -218
rect 2520 -225 2529 -222
rect 2419 -229 2463 -226
rect 2366 -245 2375 -242
rect 2419 -242 2422 -229
rect 2429 -237 2436 -234
rect 2415 -245 2422 -242
rect 2366 -278 2369 -245
rect 2419 -250 2422 -245
rect 2433 -265 2436 -237
rect 2503 -238 2506 -230
rect 2520 -234 2529 -231
rect 2520 -238 2523 -234
rect 2541 -245 2544 -211
rect 2460 -248 2544 -245
rect 2460 -252 2463 -248
rect 2528 -252 2531 -248
rect 2445 -265 2448 -260
rect 2433 -268 2448 -265
rect 2366 -281 2439 -278
rect 2366 -333 2369 -281
rect 2436 -307 2439 -281
rect 2445 -284 2448 -268
rect 2496 -265 2499 -260
rect 2457 -268 2515 -265
rect 2512 -284 2515 -268
rect 2460 -298 2463 -292
rect 2496 -298 2499 -292
rect 2528 -298 2531 -292
rect 2460 -301 2531 -298
rect 2460 -307 2463 -301
rect 2399 -318 2402 -307
rect 2436 -310 2463 -307
rect 2460 -314 2463 -310
rect 2460 -317 2531 -314
rect 2383 -321 2407 -318
rect 2460 -323 2463 -317
rect 2366 -336 2375 -333
rect 2366 -369 2369 -336
rect 2399 -369 2402 -330
rect 2496 -323 2499 -317
rect 2528 -323 2531 -317
rect 2415 -336 2422 -333
rect 2366 -372 2375 -369
rect 2366 -401 2369 -372
rect 2399 -372 2407 -369
rect 2399 -385 2402 -372
rect 2383 -388 2402 -385
rect 2419 -385 2422 -336
rect 2445 -347 2448 -331
rect 2433 -350 2448 -347
rect 2433 -376 2436 -350
rect 2445 -355 2448 -350
rect 2512 -347 2515 -331
rect 2457 -350 2515 -347
rect 2496 -355 2499 -350
rect 2429 -379 2436 -376
rect 2460 -367 2463 -363
rect 2528 -367 2531 -363
rect 2541 -367 2544 -248
rect 2460 -370 2544 -367
rect 2460 -385 2463 -370
rect 2503 -383 2506 -377
rect 2520 -381 2523 -377
rect 2419 -388 2463 -385
rect 2520 -384 2529 -381
rect 2366 -404 2375 -401
rect 2419 -401 2422 -388
rect 2429 -396 2436 -393
rect 2415 -404 2422 -401
rect 2366 -416 2369 -404
rect 2419 -409 2422 -404
rect 2366 -419 2423 -416
rect 2366 -422 2369 -419
rect 2307 -450 2414 -447
rect 2272 -462 2278 -459
rect 2275 -495 2278 -462
rect 2411 -466 2414 -450
rect 2420 -457 2423 -419
rect 2433 -424 2436 -396
rect 2503 -397 2506 -388
rect 2520 -393 2529 -390
rect 2520 -397 2523 -393
rect 2541 -404 2544 -370
rect 2549 -389 2552 82
rect 2556 -230 2559 82
rect 2563 -76 2566 82
rect 2460 -407 2544 -404
rect 2460 -411 2463 -407
rect 2528 -411 2531 -407
rect 2445 -424 2448 -419
rect 2433 -427 2448 -424
rect 2445 -443 2448 -427
rect 2496 -424 2499 -419
rect 2457 -427 2515 -424
rect 2512 -443 2515 -427
rect 2460 -457 2463 -451
rect 2496 -457 2499 -451
rect 2528 -457 2531 -451
rect 2420 -460 2531 -457
rect 2541 -466 2544 -407
rect 2411 -469 2544 -466
rect 2275 -498 2343 -495
rect 2165 -514 2189 -511
rect 2253 -514 2277 -511
rect 2064 -529 2157 -526
rect 2070 -567 2073 -529
rect 2032 -570 2040 -567
rect 2037 -583 2040 -570
rect 2064 -570 2073 -567
rect 2037 -586 2056 -583
rect 1784 -614 1787 -602
rect 1980 -614 1983 -602
rect 2017 -602 2024 -599
rect 2070 -599 2073 -570
rect 2064 -602 2073 -599
rect 2148 -567 2151 -529
rect 2181 -567 2184 -523
rect 2197 -529 2205 -526
rect 2237 -529 2245 -526
rect 2148 -570 2157 -567
rect 2148 -599 2151 -570
rect 2181 -570 2189 -567
rect 2181 -583 2184 -570
rect 2165 -586 2184 -583
rect 2148 -602 2157 -599
rect 2201 -599 2204 -529
rect 2211 -577 2219 -574
rect 2224 -577 2231 -574
rect 2211 -594 2217 -591
rect 2197 -602 2204 -599
rect 2214 -600 2217 -594
rect 2225 -594 2231 -591
rect 2225 -600 2228 -594
rect 2238 -599 2241 -529
rect 2258 -567 2261 -523
rect 2299 -526 2302 -506
rect 2340 -514 2343 -498
rect 2335 -517 2359 -514
rect 2285 -529 2302 -526
rect 2291 -567 2294 -529
rect 2253 -570 2261 -567
rect 2258 -583 2261 -570
rect 2285 -570 2294 -567
rect 2258 -586 2277 -583
rect 2017 -614 2020 -602
rect 2201 -614 2204 -602
rect 2238 -602 2245 -599
rect 2291 -599 2294 -570
rect 2320 -532 2327 -529
rect 2307 -580 2313 -577
rect 2285 -602 2294 -599
rect 2303 -597 2313 -594
rect 2238 -614 2241 -602
rect 2303 -603 2306 -597
rect 2320 -602 2323 -532
rect 2340 -570 2343 -526
rect 2379 -529 2382 -506
rect 2367 -532 2382 -529
rect 2373 -570 2376 -532
rect 2335 -573 2343 -570
rect 2340 -586 2343 -573
rect 2367 -573 2376 -570
rect 2340 -589 2359 -586
rect 2320 -605 2327 -602
rect 2373 -602 2376 -573
rect 2367 -605 2376 -602
rect 2320 -614 2323 -605
rect 1441 -615 2323 -614
rect 2411 -615 2414 -469
rect 1441 -617 2414 -615
rect 1441 -630 1444 -617
rect 2320 -618 2414 -617
rect 723 -633 1444 -630
rect 2303 -633 2306 -627
rect 956 -636 959 -633
rect 987 -636 990 -633
rect 1501 -636 2306 -633
rect 610 -643 620 -640
rect 1501 -639 1504 -636
rect 718 -642 1504 -639
rect 588 -653 605 -650
rect 538 -658 564 -655
rect 617 -661 620 -643
rect 610 -664 620 -661
rect 550 -672 553 -666
rect 572 -672 577 -664
rect 550 -675 577 -672
rect 617 -675 620 -664
rect 691 -649 806 -646
rect 560 -683 563 -675
rect 617 -678 687 -675
rect 560 -686 680 -683
rect 486 -693 673 -690
rect 444 -700 666 -697
rect 417 -707 659 -704
rect 656 -742 659 -707
rect 663 -742 666 -700
rect 670 -742 673 -693
rect 677 -742 680 -686
rect 684 -742 687 -678
rect 691 -742 694 -649
rect 811 -649 1520 -646
rect 2549 -646 2552 -394
rect 1525 -649 2552 -646
rect 698 -656 962 -653
rect 698 -742 701 -656
rect 967 -656 1759 -653
rect 2556 -653 2559 -235
rect 1764 -656 2559 -653
rect 705 -663 1112 -660
rect 705 -742 708 -663
rect 1117 -663 1992 -660
rect 2563 -660 2566 -81
rect 1997 -663 2566 -660
rect 712 -670 1268 -667
rect 712 -742 715 -670
rect 1273 -670 2213 -667
rect 2570 -667 2573 78
rect 2577 -380 2580 82
rect 2584 -221 2587 82
rect 2591 -67 2594 82
rect 2218 -670 2573 -667
rect 719 -677 823 -674
rect 719 -742 722 -677
rect 828 -677 1532 -674
rect 2577 -674 2580 -385
rect 1537 -677 2580 -674
rect 726 -684 979 -681
rect 726 -742 729 -684
rect 984 -684 1770 -681
rect 2584 -681 2587 -226
rect 1775 -684 2587 -681
rect 733 -691 1129 -688
rect 733 -742 736 -691
rect 1134 -691 2003 -688
rect 2591 -688 2594 -72
rect 2008 -691 2594 -688
rect 740 -698 1285 -695
rect 740 -742 743 -698
rect 1290 -698 2224 -695
rect 2598 -695 2601 87
rect 2229 -698 2601 -695
<< m2contact >>
rect 1050 277 1055 282
rect 1084 269 1089 274
rect 952 169 957 174
rect 1017 202 1022 207
rect 1004 172 1009 177
rect 905 137 910 142
rect 905 120 910 125
rect 751 77 756 82
rect 751 67 756 72
rect 1038 202 1043 207
rect 1135 191 1140 196
rect 1145 180 1150 185
rect 1165 195 1170 200
rect 1171 179 1176 184
rect 1368 222 1373 227
rect 1194 193 1199 198
rect 1024 135 1029 141
rect 964 119 969 124
rect 964 109 969 114
rect 924 82 929 87
rect 1163 163 1168 168
rect 1187 150 1192 155
rect 1095 105 1100 110
rect 1095 95 1100 100
rect 924 49 929 54
rect 836 26 841 31
rect 758 -8 763 -3
rect 782 -32 787 -27
rect 790 -90 795 -85
rect 807 -60 812 -55
rect 807 -70 812 -65
rect 924 28 929 33
rect 878 -85 883 -80
rect 980 23 985 28
rect 895 -55 900 -50
rect 895 -65 900 -60
rect 814 -143 819 -138
rect 795 -155 800 -150
rect 830 -162 835 -157
rect 814 -180 819 -175
rect 549 -300 554 -295
rect 534 -307 539 -302
rect 549 -334 554 -329
rect 616 -352 621 -347
rect 616 -376 621 -371
rect 549 -413 554 -408
rect 508 -420 513 -415
rect 454 -473 459 -468
rect 443 -538 448 -533
rect 513 -491 518 -486
rect 485 -548 490 -543
rect 474 -580 479 -575
rect 424 -610 429 -605
rect 443 -618 448 -613
rect 549 -447 554 -442
rect 616 -465 621 -460
rect 616 -489 621 -484
rect 549 -508 554 -503
rect 534 -528 539 -523
rect 534 -538 539 -533
rect 534 -548 539 -543
rect 549 -555 554 -550
rect 834 -235 839 -230
rect 899 -138 904 -133
rect 951 -141 956 -136
rect 918 -150 923 -145
rect 891 -174 896 -169
rect 996 23 1001 28
rect 1078 75 1083 80
rect 1292 125 1297 130
rect 1292 115 1297 120
rect 1091 -8 1096 -3
rect 1183 18 1188 23
rect 1172 13 1177 18
rect 1118 1 1123 6
rect 1071 -18 1076 -13
rect 1109 -18 1114 -13
rect 1100 -76 1105 -71
rect 1249 34 1254 39
rect 1296 34 1301 39
rect 1257 23 1262 28
rect 1321 18 1326 23
rect 1123 -46 1128 -41
rect 1123 -56 1128 -51
rect 1208 -78 1213 -73
rect 1225 -48 1230 -43
rect 1225 -58 1230 -53
rect 1126 -129 1131 -124
rect 1146 -144 1151 -139
rect 1126 -151 1131 -146
rect 834 -260 839 -255
rect 899 -262 904 -257
rect 882 -280 887 -275
rect 891 -280 896 -275
rect 845 -313 850 -308
rect 781 -338 786 -333
rect 831 -366 836 -361
rect 757 -433 762 -428
rect 809 -394 814 -389
rect 863 -428 868 -423
rect 793 -476 798 -471
rect 1020 -225 1025 -220
rect 1248 -141 1253 -136
rect 1281 -161 1286 -156
rect 1239 -169 1244 -164
rect 1311 -161 1316 -156
rect 1284 -181 1289 -176
rect 1622 348 1627 353
rect 1463 126 1468 131
rect 1679 348 1684 353
rect 1761 347 1766 352
rect 1803 347 1808 352
rect 1910 346 1915 351
rect 1949 346 1954 351
rect 1574 237 1579 242
rect 1549 211 1554 216
rect 1682 281 1687 286
rect 1694 264 1699 269
rect 1728 281 1733 286
rect 1826 283 1831 288
rect 1714 260 1719 265
rect 1838 259 1843 264
rect 1703 246 1708 251
rect 1727 246 1732 251
rect 1528 176 1533 181
rect 1637 177 1642 182
rect 1872 283 1877 288
rect 1969 284 1974 289
rect 1981 273 1986 278
rect 1858 259 1863 264
rect 2015 284 2020 289
rect 2001 274 2006 279
rect 1787 211 1792 216
rect 1766 179 1771 184
rect 1872 177 1877 182
rect 2020 214 2025 219
rect 1999 179 2004 184
rect 2108 180 2113 185
rect 2258 214 2263 219
rect 2237 182 2242 187
rect 1578 148 1583 153
rect 1504 82 1509 87
rect 1556 120 1561 125
rect 1450 46 1455 51
rect 1450 -14 1455 -9
rect 1610 86 1615 91
rect 1540 38 1545 43
rect 1701 129 1706 134
rect 1816 151 1821 156
rect 1742 85 1747 90
rect 1794 123 1799 128
rect 1688 49 1693 54
rect 1495 -56 1500 -51
rect 1514 -56 1519 -51
rect 1528 -48 1533 -43
rect 1578 -76 1583 -71
rect 1624 -87 1629 -82
rect 1022 -287 1027 -282
rect 898 -366 903 -361
rect 1034 -304 1039 -299
rect 1043 -304 1048 -299
rect 999 -313 1004 -308
rect 937 -338 942 -333
rect 987 -366 992 -361
rect 913 -433 918 -428
rect 965 -394 970 -389
rect 1019 -428 1024 -423
rect 949 -476 954 -471
rect 1050 -366 1055 -361
rect 1331 -202 1336 -197
rect 1172 -287 1177 -282
rect 1182 -307 1187 -302
rect 1191 -307 1196 -302
rect 1151 -313 1156 -308
rect 1087 -338 1092 -333
rect 1137 -366 1142 -361
rect 1063 -433 1068 -428
rect 1115 -394 1120 -389
rect 1169 -428 1174 -423
rect 739 -507 744 -502
rect 1099 -476 1104 -471
rect 1198 -366 1203 -361
rect 1271 -301 1276 -296
rect 1442 -151 1447 -146
rect 1491 -134 1496 -129
rect 1556 -104 1561 -99
rect 1504 -151 1509 -146
rect 1610 -138 1615 -133
rect 1540 -186 1545 -181
rect 1519 -214 1524 -209
rect 1557 -214 1562 -209
rect 1491 -223 1496 -218
rect 1348 -266 1353 -261
rect 1337 -293 1342 -288
rect 1234 -338 1239 -333
rect 1284 -366 1289 -361
rect 1210 -433 1215 -428
rect 1262 -394 1267 -389
rect 1316 -428 1321 -423
rect 893 -507 898 -502
rect 717 -555 722 -550
rect 702 -565 707 -560
rect 616 -572 621 -567
rect 663 -578 668 -573
rect 521 -584 526 -579
rect 504 -610 509 -605
rect 616 -594 621 -589
rect 549 -630 554 -625
rect 533 -639 538 -634
rect 485 -649 490 -644
rect 533 -649 538 -644
rect 443 -659 448 -654
rect 816 -589 821 -584
rect 1246 -476 1251 -471
rect 1046 -507 1051 -502
rect 972 -589 977 -584
rect 806 -626 811 -621
rect 823 -626 828 -621
rect 1198 -507 1203 -502
rect 1122 -589 1127 -584
rect 962 -626 967 -621
rect 979 -626 984 -621
rect 1451 -280 1456 -275
rect 1429 -308 1434 -303
rect 1501 -308 1506 -303
rect 1427 -370 1432 -365
rect 1479 -336 1484 -331
rect 1533 -370 1538 -365
rect 1463 -418 1468 -413
rect 1548 -411 1553 -406
rect 1471 -463 1476 -458
rect 1410 -507 1415 -502
rect 1364 -515 1369 -510
rect 1277 -589 1282 -584
rect 1112 -626 1117 -621
rect 1129 -626 1134 -621
rect 1688 -11 1693 -6
rect 1848 89 1853 94
rect 1778 41 1783 46
rect 1934 129 1939 134
rect 2049 151 2054 156
rect 1975 85 1980 90
rect 2027 123 2032 128
rect 1921 49 1926 54
rect 1733 -53 1738 -48
rect 1752 -53 1757 -48
rect 1766 -45 1771 -40
rect 1816 -73 1821 -68
rect 1862 -84 1867 -79
rect 1680 -148 1685 -143
rect 1729 -131 1734 -126
rect 1794 -101 1799 -96
rect 1742 -148 1747 -143
rect 1848 -135 1853 -130
rect 1778 -183 1783 -178
rect 1757 -211 1762 -206
rect 1795 -211 1800 -206
rect 1729 -220 1734 -215
rect 1590 -308 1595 -303
rect 1689 -277 1694 -272
rect 1667 -305 1672 -300
rect 1739 -305 1744 -300
rect 1665 -371 1670 -366
rect 1717 -333 1722 -328
rect 1771 -367 1776 -362
rect 1701 -415 1706 -410
rect 1786 -415 1791 -410
rect 1709 -463 1714 -458
rect 1635 -506 1640 -501
rect 1364 -538 1369 -533
rect 1364 -565 1369 -560
rect 1526 -579 1531 -574
rect 1921 -11 1926 -6
rect 2081 89 2086 94
rect 2011 41 2016 46
rect 2172 132 2177 137
rect 2287 154 2292 159
rect 2399 160 2404 165
rect 2213 88 2218 93
rect 2265 126 2270 131
rect 2159 52 2164 57
rect 1966 -53 1971 -48
rect 1985 -53 1990 -48
rect 1999 -45 2004 -40
rect 2049 -73 2054 -68
rect 2095 -84 2100 -79
rect 1913 -148 1918 -143
rect 1962 -131 1967 -126
rect 2027 -101 2032 -96
rect 1975 -148 1980 -143
rect 2081 -135 2086 -130
rect 2011 -183 2016 -178
rect 1990 -211 1995 -206
rect 2028 -211 2033 -206
rect 1962 -220 1967 -215
rect 1828 -305 1833 -300
rect 1922 -277 1927 -272
rect 1900 -305 1905 -300
rect 1972 -305 1977 -300
rect 1898 -372 1903 -367
rect 1950 -333 1955 -328
rect 2004 -367 2009 -362
rect 1934 -415 1939 -410
rect 2019 -414 2024 -409
rect 1942 -463 1947 -458
rect 1861 -506 1866 -501
rect 1268 -625 1273 -620
rect 1285 -625 1290 -620
rect 1520 -606 1525 -601
rect 1532 -606 1537 -601
rect 1765 -578 1770 -573
rect 2159 -8 2164 -3
rect 2319 92 2324 97
rect 2249 44 2254 49
rect 2503 83 2508 88
rect 2530 87 2535 92
rect 2530 78 2535 83
rect 2597 87 2602 92
rect 2204 -50 2209 -45
rect 2223 -50 2228 -45
rect 2399 7 2404 12
rect 2237 -42 2242 -37
rect 2287 -70 2292 -65
rect 2333 -81 2338 -76
rect 2151 -145 2156 -140
rect 2200 -128 2205 -123
rect 2265 -98 2270 -93
rect 2213 -145 2218 -140
rect 2319 -132 2324 -127
rect 2249 -180 2254 -175
rect 2228 -208 2233 -203
rect 2266 -208 2271 -203
rect 2200 -217 2205 -212
rect 2061 -305 2066 -300
rect 2160 -274 2165 -269
rect 2138 -302 2143 -297
rect 2210 -302 2215 -297
rect 2136 -368 2141 -363
rect 2188 -330 2193 -325
rect 2242 -364 2247 -359
rect 2172 -412 2177 -407
rect 2104 -506 2109 -501
rect 1759 -605 1764 -600
rect 1770 -605 1775 -600
rect 1998 -578 2003 -573
rect 2197 -455 2202 -450
rect 2267 -463 2272 -458
rect 2503 -75 2508 -70
rect 2530 -72 2535 -67
rect 2530 -81 2535 -76
rect 2398 -147 2403 -142
rect 2299 -302 2304 -297
rect 2502 -230 2507 -225
rect 2529 -226 2534 -221
rect 2529 -235 2534 -230
rect 2398 -307 2403 -302
rect 2502 -388 2507 -383
rect 2529 -385 2534 -380
rect 2365 -427 2370 -422
rect 2529 -394 2534 -389
rect 2569 78 2574 83
rect 2562 -81 2567 -76
rect 2555 -235 2560 -230
rect 2548 -394 2553 -389
rect 2298 -506 2303 -501
rect 1992 -605 1997 -600
rect 2003 -605 2008 -600
rect 2219 -578 2224 -573
rect 2378 -506 2383 -501
rect 2213 -605 2218 -600
rect 2224 -605 2229 -600
rect 2302 -581 2307 -576
rect 2302 -608 2307 -603
rect 2302 -627 2307 -622
rect 713 -643 718 -638
rect 533 -659 538 -654
rect 549 -666 554 -661
rect 412 -708 417 -703
rect 806 -650 811 -645
rect 1520 -650 1525 -645
rect 962 -657 967 -652
rect 1759 -657 1764 -652
rect 1112 -664 1117 -659
rect 1992 -664 1997 -659
rect 1268 -671 1273 -666
rect 2213 -671 2218 -666
rect 2590 -72 2595 -67
rect 2583 -226 2588 -221
rect 2576 -385 2581 -380
rect 823 -678 828 -673
rect 1532 -678 1537 -673
rect 979 -685 984 -680
rect 1770 -685 1775 -680
rect 1129 -692 1134 -687
rect 2003 -692 2008 -687
rect 1285 -699 1290 -694
rect 2224 -699 2229 -694
<< metal2 >>
rect 1627 349 1679 352
rect 1766 348 1803 351
rect 1915 347 1949 350
rect 1687 282 1728 285
rect 1831 284 1872 287
rect 1974 285 2015 288
rect 1055 278 1541 281
rect 1538 277 1541 278
rect 1538 274 1981 277
rect 1096 273 1500 274
rect 1089 271 1500 273
rect 1089 270 1099 271
rect 1497 268 1500 271
rect 1497 265 1694 268
rect 1566 247 1703 250
rect 1566 232 1569 247
rect 1715 240 1718 260
rect 1839 250 1842 259
rect 1732 247 1842 250
rect 1859 247 1862 259
rect 2002 254 2005 274
rect 2002 251 2371 254
rect 1859 244 2364 247
rect 1715 237 2357 240
rect 1535 229 1569 232
rect 1575 233 1578 237
rect 1575 230 2350 233
rect 1535 226 1538 229
rect 1373 223 1538 226
rect 1812 224 2262 226
rect 1550 223 2262 224
rect 1550 221 1815 223
rect 1550 216 1553 221
rect 1788 216 1791 221
rect 2021 219 2024 223
rect 2259 219 2262 223
rect 1022 203 1038 206
rect 917 192 1135 195
rect 906 125 909 137
rect 735 78 751 81
rect 735 -151 738 78
rect 917 76 920 192
rect 1170 196 1183 199
rect 925 181 1145 184
rect 925 87 928 181
rect 1009 174 1043 177
rect 953 140 956 169
rect 1040 167 1043 174
rect 1040 164 1163 167
rect 953 136 1024 140
rect 948 120 964 123
rect 837 73 920 76
rect 742 68 751 71
rect 742 63 745 68
rect 742 60 751 63
rect 748 -104 751 60
rect 837 31 840 73
rect 948 66 951 120
rect 955 110 964 113
rect 955 105 958 110
rect 1079 106 1095 109
rect 955 102 964 105
rect 879 63 951 66
rect 759 -28 762 -8
rect 759 -31 782 -28
rect 879 -51 882 63
rect 925 33 928 49
rect 879 -54 895 -51
rect 791 -59 807 -56
rect 791 -85 794 -59
rect 798 -69 807 -66
rect 798 -74 801 -69
rect 798 -77 807 -74
rect 804 -104 807 -77
rect 879 -80 882 -54
rect 886 -64 895 -61
rect 886 -69 889 -64
rect 886 -72 895 -69
rect 748 -108 807 -104
rect 735 -154 795 -151
rect 804 -265 807 -108
rect 815 -175 818 -143
rect 831 -166 834 -162
rect 831 -169 857 -166
rect 892 -169 895 -72
rect 835 -255 838 -235
rect 804 -268 815 -265
rect 812 -300 815 -268
rect 854 -266 857 -169
rect 854 -269 886 -266
rect 883 -275 886 -269
rect 892 -275 895 -174
rect 900 -257 903 -138
rect 911 -140 951 -137
rect 911 -221 914 -140
rect 919 -161 922 -150
rect 961 -161 964 102
rect 1079 80 1082 106
rect 1086 96 1095 99
rect 1086 91 1089 96
rect 1086 88 1095 91
rect 985 24 996 27
rect 1092 -3 1095 88
rect 1172 18 1175 179
rect 1180 64 1183 196
rect 1195 188 1198 193
rect 1188 185 1198 188
rect 1188 155 1191 185
rect 1529 152 1532 176
rect 1498 149 1532 152
rect 1498 138 1501 149
rect 1529 148 1532 149
rect 1583 149 1622 152
rect 1529 145 1560 148
rect 1496 134 1501 138
rect 1464 131 1499 134
rect 1276 126 1292 129
rect 1180 61 1261 64
rect 1217 35 1249 38
rect 1217 22 1220 35
rect 1258 28 1261 61
rect 1188 19 1220 22
rect 1276 15 1279 126
rect 1557 125 1560 145
rect 1283 116 1292 119
rect 1283 111 1286 116
rect 1283 108 1292 111
rect 1209 12 1279 15
rect 1289 15 1292 108
rect 1607 87 1610 149
rect 1505 77 1508 82
rect 1611 79 1614 86
rect 1505 74 1522 77
rect 1519 50 1522 74
rect 1599 76 1614 79
rect 1599 50 1602 76
rect 1519 47 1602 50
rect 1297 22 1300 34
rect 1297 19 1321 22
rect 1289 12 1299 15
rect 1076 -17 1109 -14
rect 1119 -34 1122 1
rect 1093 -37 1122 -34
rect 1093 -160 1096 -37
rect 1101 -45 1123 -42
rect 1101 -71 1104 -45
rect 1209 -44 1212 12
rect 1209 -47 1225 -44
rect 1114 -55 1123 -52
rect 1114 -160 1117 -55
rect 1209 -73 1212 -47
rect 1216 -57 1225 -54
rect 1216 -62 1219 -57
rect 1216 -65 1225 -62
rect 1127 -146 1130 -129
rect 1147 -152 1150 -144
rect 1147 -155 1186 -152
rect 919 -165 1038 -161
rect 911 -224 1020 -221
rect 413 -306 534 -303
rect 413 -416 416 -306
rect 550 -329 553 -300
rect 812 -303 857 -300
rect 854 -309 857 -303
rect 850 -312 919 -309
rect 617 -371 620 -352
rect 782 -362 785 -338
rect 729 -365 785 -362
rect 413 -419 508 -416
rect 413 -524 416 -419
rect 550 -442 553 -413
rect 455 -464 616 -461
rect 455 -468 458 -464
rect 617 -477 620 -465
rect 729 -477 732 -365
rect 782 -366 785 -365
rect 836 -365 898 -362
rect 782 -369 813 -366
rect 810 -389 813 -369
rect 860 -427 863 -365
rect 916 -362 919 -312
rect 1023 -309 1026 -287
rect 1035 -299 1038 -165
rect 1087 -163 1117 -160
rect 1087 -257 1090 -163
rect 1044 -260 1090 -257
rect 1044 -299 1047 -260
rect 1004 -312 1069 -309
rect 938 -362 941 -338
rect 916 -365 941 -362
rect 938 -366 941 -365
rect 992 -365 1050 -362
rect 938 -369 969 -366
rect 966 -389 969 -369
rect 1016 -427 1019 -365
rect 1066 -362 1069 -312
rect 1156 -311 1163 -309
rect 1173 -311 1176 -287
rect 1183 -302 1186 -155
rect 1222 -165 1225 -65
rect 1249 -145 1252 -141
rect 1295 -145 1299 12
rect 1451 -2 1454 46
rect 1541 43 1544 47
rect 1451 -5 1465 -2
rect 1451 -9 1454 -5
rect 1462 -87 1465 -5
rect 1500 -55 1514 -52
rect 1529 -72 1532 -48
rect 1507 -75 1532 -72
rect 1507 -82 1511 -75
rect 1529 -76 1532 -75
rect 1598 -72 1601 47
rect 1583 -75 1628 -72
rect 1529 -79 1560 -76
rect 1500 -85 1511 -82
rect 1500 -87 1504 -85
rect 1249 -149 1299 -145
rect 1453 -90 1504 -87
rect 1222 -168 1239 -165
rect 1222 -263 1225 -168
rect 1249 -182 1252 -149
rect 1453 -147 1456 -90
rect 1557 -99 1560 -79
rect 1447 -150 1456 -147
rect 1286 -160 1311 -157
rect 1289 -180 1335 -177
rect 1248 -185 1252 -182
rect 1192 -266 1225 -263
rect 1192 -302 1195 -266
rect 1249 -272 1252 -185
rect 1332 -197 1335 -180
rect 1492 -218 1495 -134
rect 1607 -137 1610 -75
rect 1625 -82 1628 -75
rect 1611 -145 1614 -138
rect 1599 -148 1614 -145
rect 1505 -155 1508 -151
rect 1505 -158 1522 -155
rect 1519 -174 1522 -158
rect 1599 -174 1602 -148
rect 1519 -177 1602 -174
rect 1541 -181 1544 -177
rect 1524 -213 1557 -210
rect 1323 -265 1348 -262
rect 1249 -275 1264 -272
rect 1261 -289 1264 -275
rect 1323 -281 1326 -265
rect 1323 -284 1351 -281
rect 1261 -292 1337 -289
rect 1276 -300 1297 -297
rect 1348 -298 1351 -284
rect 1156 -312 1216 -311
rect 1160 -314 1216 -312
rect 1088 -362 1091 -338
rect 1066 -365 1091 -362
rect 1088 -366 1091 -365
rect 1142 -365 1198 -362
rect 1088 -369 1119 -366
rect 1116 -389 1119 -369
rect 1166 -427 1169 -365
rect 1213 -362 1216 -314
rect 1235 -362 1238 -338
rect 1213 -365 1238 -362
rect 1235 -366 1238 -365
rect 1294 -362 1297 -300
rect 1326 -301 1351 -298
rect 1326 -362 1329 -301
rect 1452 -304 1455 -280
rect 1434 -307 1455 -304
rect 1452 -308 1455 -307
rect 1506 -307 1590 -304
rect 1452 -311 1483 -308
rect 1480 -331 1483 -311
rect 1289 -365 1348 -362
rect 1235 -369 1266 -366
rect 1263 -389 1266 -369
rect 1313 -427 1316 -365
rect 1345 -389 1348 -365
rect 1530 -369 1533 -307
rect 1428 -379 1431 -370
rect 1534 -377 1537 -370
rect 1428 -382 1445 -379
rect 1442 -389 1445 -382
rect 1345 -392 1445 -389
rect 1442 -406 1445 -392
rect 1522 -380 1537 -377
rect 1522 -406 1525 -380
rect 1442 -409 1525 -406
rect 1464 -413 1467 -409
rect 1549 -415 1552 -411
rect 1638 -415 1641 177
rect 1767 155 1770 179
rect 1736 152 1770 155
rect 1736 141 1739 152
rect 1767 151 1770 152
rect 1821 152 1860 155
rect 1767 148 1798 151
rect 1734 137 1739 141
rect 1702 134 1737 137
rect 1795 128 1798 148
rect 1845 90 1848 152
rect 1743 80 1746 85
rect 1849 82 1852 89
rect 1743 77 1760 80
rect 1757 53 1760 77
rect 1837 79 1852 82
rect 1837 53 1840 79
rect 1757 50 1840 53
rect 1689 1 1692 49
rect 1779 46 1782 50
rect 1689 -2 1703 1
rect 1689 -6 1692 -2
rect 1700 -84 1703 -2
rect 1738 -52 1752 -49
rect 1767 -69 1770 -45
rect 1745 -72 1770 -69
rect 1745 -79 1749 -72
rect 1767 -73 1770 -72
rect 1836 -69 1839 50
rect 1821 -72 1866 -69
rect 1767 -76 1798 -73
rect 1738 -82 1749 -79
rect 1738 -84 1742 -82
rect 1691 -87 1742 -84
rect 1691 -144 1694 -87
rect 1795 -96 1798 -76
rect 1685 -147 1694 -144
rect 1730 -215 1733 -131
rect 1845 -134 1848 -72
rect 1863 -79 1866 -72
rect 1849 -142 1852 -135
rect 1837 -145 1852 -142
rect 1743 -152 1746 -148
rect 1743 -155 1760 -152
rect 1757 -171 1760 -155
rect 1837 -171 1840 -145
rect 1757 -174 1840 -171
rect 1779 -178 1782 -174
rect 1762 -210 1795 -207
rect 1690 -301 1693 -277
rect 1672 -304 1693 -301
rect 1690 -305 1693 -304
rect 1744 -304 1828 -301
rect 1690 -308 1721 -305
rect 1718 -328 1721 -308
rect 1768 -366 1771 -304
rect 1666 -376 1669 -371
rect 1772 -374 1775 -367
rect 1666 -379 1683 -376
rect 1680 -403 1683 -379
rect 1760 -377 1775 -374
rect 1760 -403 1763 -377
rect 1680 -406 1763 -403
rect 1702 -410 1705 -406
rect 1549 -418 1641 -415
rect 1787 -419 1790 -415
rect 1873 -419 1876 177
rect 2000 155 2003 179
rect 1969 152 2003 155
rect 1969 141 1972 152
rect 2000 151 2003 152
rect 2054 152 2093 155
rect 2000 148 2031 151
rect 1967 137 1972 141
rect 1935 134 1970 137
rect 2028 128 2031 148
rect 2078 90 2081 152
rect 1976 80 1979 85
rect 2082 82 2085 89
rect 1976 77 1993 80
rect 1990 53 1993 77
rect 2070 79 2085 82
rect 2070 53 2073 79
rect 1990 50 2073 53
rect 1922 1 1925 49
rect 2012 46 2015 50
rect 1922 -2 1936 1
rect 1922 -6 1925 -2
rect 1933 -84 1936 -2
rect 1971 -52 1985 -49
rect 2000 -69 2003 -45
rect 1978 -72 2003 -69
rect 1978 -79 1982 -72
rect 2000 -73 2003 -72
rect 2069 -69 2072 50
rect 2054 -72 2099 -69
rect 2000 -76 2031 -73
rect 1971 -82 1982 -79
rect 1971 -84 1975 -82
rect 1924 -87 1975 -84
rect 1924 -144 1927 -87
rect 2028 -96 2031 -76
rect 1918 -147 1927 -144
rect 1963 -215 1966 -131
rect 2078 -134 2081 -72
rect 2096 -79 2099 -72
rect 2082 -142 2085 -135
rect 2070 -145 2085 -142
rect 1976 -152 1979 -148
rect 1976 -155 1993 -152
rect 1990 -171 1993 -155
rect 2070 -171 2073 -145
rect 1990 -174 2073 -171
rect 2012 -178 2015 -174
rect 1995 -210 2028 -207
rect 1923 -301 1926 -277
rect 1905 -304 1926 -301
rect 1923 -305 1926 -304
rect 1977 -304 2061 -301
rect 1923 -308 1954 -305
rect 1951 -328 1954 -308
rect 2001 -366 2004 -304
rect 1899 -376 1902 -372
rect 2005 -374 2008 -367
rect 1899 -379 1916 -376
rect 1913 -403 1916 -379
rect 1993 -377 2008 -374
rect 1993 -403 1996 -377
rect 1913 -406 1996 -403
rect 1935 -410 1938 -406
rect 1787 -422 1876 -419
rect 2020 -418 2023 -414
rect 2109 -418 2112 180
rect 2238 158 2241 182
rect 2207 155 2241 158
rect 2207 144 2210 155
rect 2238 154 2241 155
rect 2292 155 2331 158
rect 2238 151 2269 154
rect 2205 140 2210 144
rect 2173 137 2208 140
rect 2266 131 2269 151
rect 2316 93 2319 155
rect 2214 83 2217 88
rect 2320 85 2323 92
rect 2214 80 2231 83
rect 2228 56 2231 80
rect 2308 82 2323 85
rect 2308 56 2311 82
rect 2228 53 2311 56
rect 2160 4 2163 52
rect 2250 49 2253 53
rect 2160 1 2174 4
rect 2160 -3 2163 1
rect 2171 -81 2174 1
rect 2209 -49 2223 -46
rect 2238 -66 2241 -42
rect 2216 -69 2241 -66
rect 2216 -76 2220 -69
rect 2238 -70 2241 -69
rect 2307 -66 2310 53
rect 2292 -69 2337 -66
rect 2238 -73 2269 -70
rect 2209 -79 2220 -76
rect 2209 -81 2213 -79
rect 2162 -84 2213 -81
rect 2162 -141 2165 -84
rect 2266 -93 2269 -73
rect 2156 -144 2165 -141
rect 2201 -212 2204 -128
rect 2316 -131 2319 -69
rect 2334 -76 2337 -69
rect 2320 -139 2323 -132
rect 2308 -142 2323 -139
rect 2214 -149 2217 -145
rect 2214 -152 2231 -149
rect 2228 -168 2231 -152
rect 2308 -168 2311 -142
rect 2228 -171 2311 -168
rect 2250 -175 2253 -171
rect 2233 -207 2266 -204
rect 2161 -298 2164 -274
rect 2143 -301 2164 -298
rect 2161 -302 2164 -301
rect 2215 -301 2299 -298
rect 2161 -305 2192 -302
rect 2189 -325 2192 -305
rect 2239 -363 2242 -301
rect 2347 -303 2350 230
rect 2354 -143 2357 237
rect 2361 11 2364 244
rect 2368 183 2371 251
rect 2368 180 2403 183
rect 2400 165 2403 180
rect 2480 84 2503 87
rect 2361 8 2399 11
rect 2480 -71 2483 84
rect 2535 88 2597 91
rect 2602 88 2603 91
rect 2535 79 2569 82
rect 2574 79 2603 82
rect 2480 -74 2503 -71
rect 2354 -146 2398 -143
rect 2480 -226 2483 -74
rect 2535 -71 2590 -68
rect 2595 -71 2603 -68
rect 2535 -80 2562 -77
rect 2567 -80 2603 -77
rect 2480 -229 2502 -226
rect 2347 -306 2398 -303
rect 2137 -373 2140 -368
rect 2243 -371 2246 -364
rect 2137 -376 2154 -373
rect 2151 -400 2154 -376
rect 2231 -374 2246 -371
rect 2231 -400 2234 -374
rect 2151 -403 2234 -400
rect 2480 -384 2483 -229
rect 2534 -225 2583 -222
rect 2588 -225 2603 -222
rect 2534 -234 2555 -231
rect 2560 -234 2603 -231
rect 2480 -387 2502 -384
rect 2173 -407 2176 -403
rect 2020 -421 2112 -418
rect 758 -437 761 -433
rect 864 -435 867 -428
rect 758 -440 775 -437
rect 772 -464 775 -440
rect 852 -438 867 -435
rect 914 -437 917 -433
rect 1020 -435 1023 -428
rect 852 -464 855 -438
rect 914 -440 931 -437
rect 772 -467 855 -464
rect 928 -464 931 -440
rect 1008 -438 1023 -435
rect 1064 -437 1067 -433
rect 1170 -435 1173 -428
rect 1008 -464 1011 -438
rect 1064 -440 1081 -437
rect 928 -467 1011 -464
rect 1078 -464 1081 -440
rect 1158 -438 1173 -435
rect 1211 -437 1214 -433
rect 1317 -435 1320 -428
rect 1158 -464 1161 -438
rect 1211 -440 1228 -437
rect 1078 -467 1161 -464
rect 1225 -464 1228 -440
rect 1305 -438 1320 -435
rect 1305 -464 1308 -438
rect 1476 -462 1709 -459
rect 1714 -462 1942 -459
rect 2198 -459 2201 -455
rect 1947 -462 2267 -459
rect 1225 -467 1308 -464
rect 794 -471 797 -467
rect 950 -471 953 -467
rect 1100 -471 1103 -467
rect 1247 -471 1250 -467
rect 617 -480 732 -477
rect 617 -484 620 -480
rect 518 -490 535 -487
rect 532 -513 535 -490
rect 729 -503 732 -480
rect 729 -506 739 -503
rect 744 -506 893 -503
rect 898 -506 1046 -503
rect 1051 -506 1198 -503
rect 1203 -506 1410 -503
rect 1616 -503 1635 -502
rect 1415 -505 1635 -503
rect 1415 -506 1620 -505
rect 1640 -505 1861 -502
rect 1866 -505 2104 -502
rect 2109 -505 2298 -502
rect 2366 -502 2369 -427
rect 2303 -505 2378 -502
rect 2383 -505 2384 -502
rect 550 -513 553 -508
rect 532 -516 553 -513
rect 413 -527 534 -524
rect 413 -635 416 -527
rect 448 -537 534 -534
rect 490 -547 534 -544
rect 550 -550 553 -516
rect 1365 -533 1368 -515
rect 2480 -542 2483 -387
rect 2534 -384 2576 -381
rect 2581 -384 2603 -381
rect 2534 -393 2548 -390
rect 2553 -393 2603 -390
rect 664 -545 2483 -542
rect 475 -571 616 -568
rect 475 -575 478 -571
rect 429 -609 504 -606
rect 522 -614 525 -584
rect 617 -589 620 -572
rect 664 -573 667 -545
rect 722 -554 2306 -551
rect 707 -564 1364 -561
rect 817 -584 820 -564
rect 973 -584 976 -564
rect 1123 -584 1126 -564
rect 1278 -584 1281 -564
rect 1527 -574 1530 -554
rect 1766 -573 1769 -554
rect 1999 -573 2002 -554
rect 2220 -573 2223 -554
rect 2303 -576 2306 -554
rect 448 -617 525 -614
rect 522 -620 717 -617
rect 413 -638 533 -635
rect 413 -703 416 -638
rect 490 -648 533 -645
rect 448 -658 533 -655
rect 550 -661 553 -630
rect 714 -638 717 -620
rect 807 -645 810 -626
rect 807 -700 810 -650
rect 824 -673 827 -626
rect 963 -652 966 -626
rect 824 -700 827 -678
rect 963 -700 966 -657
rect 980 -680 983 -626
rect 1113 -659 1116 -626
rect 980 -700 983 -685
rect 1113 -700 1116 -664
rect 1130 -687 1133 -626
rect 1269 -666 1272 -625
rect 1130 -700 1133 -692
rect 1269 -700 1272 -671
rect 1286 -694 1289 -625
rect 1521 -645 1524 -606
rect 1286 -700 1289 -699
rect 1521 -700 1524 -650
rect 1533 -673 1536 -606
rect 1760 -652 1763 -605
rect 1533 -700 1536 -678
rect 1760 -700 1763 -657
rect 1771 -680 1774 -605
rect 1993 -659 1996 -605
rect 1771 -700 1774 -685
rect 1993 -700 1996 -664
rect 2004 -687 2007 -605
rect 2214 -666 2217 -605
rect 2004 -700 2007 -692
rect 2214 -700 2217 -671
rect 2225 -694 2228 -605
rect 2303 -622 2306 -608
rect 2225 -700 2228 -699
<< labels >>
rlabel metal1 2400 -308 2401 -307 1 YA3
rlabel metal1 2400 -149 2401 -148 1 YA2
rlabel metal1 2401 5 2402 6 1 YA1
rlabel metal1 741 -741 742 -740 1 A0
rlabel metal1 734 -741 735 -740 1 A1
rlabel metal1 727 -741 728 -740 1 A2
rlabel metal1 720 -741 721 -740 1 A3
rlabel metal1 713 -741 714 -740 1 B0
rlabel metal1 706 -741 707 -740 1 B1
rlabel metal1 699 -741 700 -740 1 B2
rlabel metal1 692 -741 693 -740 1 B3
rlabel metal1 685 -741 686 -740 1 VDD
rlabel metal1 678 -741 679 -740 1 GND
rlabel metal1 671 -741 672 -740 1 S1
rlabel metal1 664 -741 665 -740 1 S0
rlabel metal1 657 -741 658 -740 1 E
rlabel metal1 2401 159 2402 160 1 YA0
rlabel metal1 1086 282 1087 284 3 L
rlabel metal1 1052 292 1053 294 3 G
rlabel metal1 1523 257 1524 259 1 SA3
rlabel metal1 1761 253 1762 255 1 SA2
rlabel metal1 1994 251 1995 253 1 SA1
rlabel metal1 2232 257 2233 259 1 SA0
rlabel metal1 1370 229 1371 231 1 EQUAL
rlabel metal1 1472 424 1473 426 5 C
rlabel metal1 1486 424 1487 426 1 Y2
rlabel metal1 1479 424 1480 426 5 Y3
rlabel metal1 1493 424 1494 426 5 Y1
rlabel metal1 1500 424 1501 426 1 Y0
<< end >>
