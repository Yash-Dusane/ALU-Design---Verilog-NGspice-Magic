*ALU CIRCUIT 

.include TSMC_180nm.txt
.include GATES.sub
.include 2to4DECODER.sub

.include ENABLE.sub
.include 4bADDERSUB.sub
.include 4bAND.sub
.include 4bCOMPARATOR.sub

.param SUPPLY = 1.8
.param ⋋ = 0.18u

.param wn1 = {10*⋋}
.param wn2 = {10*⋋}
.param ln1 = {2*⋋}
.param ln2 = {2*⋋}

.param wp1 = wn1
.param wp2 = wn1
.param lp1 = {⋋}
.param lp2 = {⋋}

.global GND

Vdd VDD GND 'SUPPLY'

Ve E GND PULSE(0 1.8 20ns 10ps 10ps 180ns 200ns)

VS0 S1 GND PULSE(0 1.8 400ns 10ps 10ps 400ns 800ns)
VS1 S0 GND PULSE(0 1.8 200ns 10ps 10ps 200ns 400ns)

Va0 A0 GND PULSE(0 1.8 20ns 10ps 10ps 20ns 60ns)
Va1 A1 GND PULSE(0 1.8 20ns 10ps 10ps 20ns 40ns)
Va2 A2 GND PULSE(0 1.8 0ns 10ps 10ps 20ns 60ns)
Va3 A3 GND PULSE(0 1.8 0ns 10ps 10ps 20ns 40ns)

Vb0 B0 GND PULSE(0 1.8 40ns 10ps 10ps 40ns 80ns)
Vb1 B1 GND PULSE(0 1.8 0ns 10ps 10ps 20ns 60ns)
Vb2 B2 GND PULSE(0 1.8 0ns 10ps 10ps 40ns 80ns)
Vb3 B3 GND PULSE(0 1.8 20ns 10ps 10ps 40ns 60ns)

Xf E S0 S1 A0 A1 A2 A3 B0 B1 B2 B3 Y0 Y1 Y2 Y3 YC VDD GND 2to4DECODER

C0 Y0 GND 10f
C1 Y1 GND 10f
C2 Y2 GND 10f
C3 Y3 GND 10f
CC YC GND 10f

.tran 1ns 800ns

.control
run
set color0 = rgb:f/f/f
set color1 = black
plot v(E)-10 v(S0)-6 v(S1)-4 v(A0) v(A1)+2 v(A2)+4 v(A3)+6 v(B0)+10 v(B1)+12 v(B2)+14 v(B3)+16 v(Y0)+20 v(Y1)+22 v(Y2)+24 v(Y3)+26 v(YC)+28 
hardcopy image.ps v(E)-10 v(S0)-6 v(S1)-4 v(A0) v(A1)+2 v(A2)+4 v(A3)+6 v(B0)+10 v(B1)+12 v(B2)+14 v(B3)+16 v(Y0)+20 v(Y1)+22 v(Y2)+24 v(Y3)+26 v(YC)+28
.endc
.end

